library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity top is
  Port ( MCLK1 : in  STD_LOGIC;
         RS_TX : out  STD_LOGIC);
end top;

architecture fpu2 of top is

   component clock
    port (
          CLKIN_IN        : in    std_logic; 
          RST_IN          : in    std_logic; 
          CLKFX_OUT       : out   std_logic; 
          CLKIN_IBUFG_OUT : out   std_logic; 
          CLK0_OUT        : out   std_logic; 
          LOCKED_OUT      : out   std_logic);
  end component;

  signal clk: std_logic;
  type input_rom is array(0 to 199) of std_logic_vector(31 downto 0);
  type output_rom is array(0 to 99) of std_logic_vector(31 downto 0);

  constant input_data: input_rom :=(
    "11000000111100111001001010101101",
    "11101100011010101101101101110000",
    "00001111110010110100011110000000",
    "10101100011000011011111100100001",
    "10000010101010111100000000011111",
    "00111100100110010111101010011010",
    "01011110001101110101001011000011",
    "00101000011001011110010100010010",
    "11010001011111011001001011010100",
    "10110110011001000010101010100001",
    "11010110000000100101111100111111",
    "10011111000111011000001111100001",
    "10111111011110110110010000011010",
    "11101010100000001001101011000011",
    "11000010001010000011011000100111",
    "01010001000101001110110000001000",
    "10100010011011001100111011010110",
    "10100100001101000100000010100100",
    "11100000110000100101101100100000",
    "11011000001111110000000100011011",
    "11101011100110110011010100010010",
    "10011011010011111011010111110111",
    "00000110000011000010011101000100",
    "00111011001111000011001111001001",
    "11010111111111101111000101001001",
    "10110000101001011101010011010001",
    "10101100000100000000110000100011",
    "00001011000010000011000011110111",
    "11001100010001110111001111111001",
    "10111110000000010101100101111001",
    "10010100101101010011100010000101",
    "00000101101110111111101000001111",
    "10101010101101000101011101101100",
    "10000011100110111111110100000011",
    "00001001000010111010110100001101",
    "01111100000101010010111001111001",
    "11101100011110101010110111011000",
    "01010100010111110111001101000010",
    "01111000111111011000100010111111",
    "10001110101100001000001000110010",
    "00000101110011100111000101100000",
    "01110011010111000011101001111010",
    "10110111100011111001101011011101",
    "01101011011001001001110010000110",
    "11110000111001101100101111100000",
    "01010111100111101011111001000011",
    "01001100111101000110000000000111",
    "11011101110101001011001101100101",
    "00100111110000100000111100010010",
    "11010101100110000010001011000110",
    "10001101001010100011111010101110",
    "10100001001001110000011100101110",
    "01011111110011000101001001101101",
    "10010100001010101010110010011111",
    "10001010011100110001010101001111",
    "01100001111010100111101000111100",
    "01001111110101000011001100100101",
    "00010001010111111110011011000001",
    "10000111111010000101011111110100",
    "01010000110001011001011010110110",
    "00101010111000000110110100011100",
    "11000000011111010100111011110111",
    "10101111111000010000101000000000",
    "10001111110001000011000001011001",
    "01000010101110001011101000110110",
    "11010100011101011101111001000010",
    "00101110000001111011010100111100",
    "00011111100001011111101111100000",
    "10111100010111010110101000100000",
    "00011100001010010111100100011010",
    "00001000110111100011000101101100",
    "00000001000100101101111101110011",
    "10110011111010010000001010110000",
    "00100100011011100001111100110000",
    "00111110101101101011001111010100",
    "10110111111101001111001001101111",
    "00001110100110001010101010010011",
    "00110001011110011011100010110010",
    "10111001110001010101000001011110",
    "01110001111010100011000100000100",
    "01010101011100100110011010001000",
    "01000111010110000010001010100101",
    "11011001100110010011000011111011",
    "00111110100011000110110100111111",
    "10011110101110000100101111111010",
    "10010011010010000100101100000100",
    "10111100111011111111000000010001",
    "10111111000011010100110101000110",
    "10010100100111101010010110011111",
    "10000011111110100010011001111110",
    "01100101000010111010010111010100",
    "00111000100101010000011001000011",
    "10011010100010111101011111101010",
    "10001100111001011000011010010100",
    "01000101101000010010011001111100",
    "11011001001101101011001010111010",
    "00110101101101000100000001011000",
    "00011010110110100101010010100101",
    "10001100001110110110101001110101",
    "01100011001100100000111100000100",
    "10011100111010011000011100000111",
    "00000001011100111101001111001100",
    "10101100000000100101101010001100",
    "10101000110100100111111010001111",
    "10011000011010011001010101111110",
    "01000001110110011100001000100001",
    "00100101010100111100100110010011",
    "10111001100011111100100101100101",
    "11001010110110000101000000011101",
    "01111101010100011110000011111101",
    "10001000110011111001111001110010",
    "00100000111000110101110000110111",
    "10011101000100001001111001010011",
    "11011100001100101000111011000011",
    "01001000010100110111000001110110",
    "10100111000100011110011000111010",
    "01100011100010110010111010110001",
    "01001110101101001010100010110111",
    "11001000100110101101110010011110",
    "10000000011001110000110001111001",
    "11101000101010110011110001001010",
    "10101110100001101111111110000100",
    "10100110100101011000001101010000",
    "10011101000101100000101111100111",
    "01011010100110111000001100111111",
    "11011011100010000100110001001100",
    "11001100101100111110011000100010",
    "11011001101010010101000111001110",
    "11111111010101011100110111000000",
    "11001110001110111001111101110011",
    "00111100100010010110000110100110",
    "01010101101111111101100110111011",
    "10110100010000111000110110000011",
    "01000001001101111000001101011010",
    "01011100000000111000011100010001",
    "00110110010000100010010110000110",
    "11110011110000100000010100110011",
    "01100110110000001000001001000001",
    "11010111000000001001010111110011",
    "10111100001110001010011101001001",
    "11101000100000011011101011010000",
    "00110111011101100000010000010110",
    "00111011010110011111100001001001",
    "11010011110000100110101011101100",
    "11010000101011001000110100010110",
    "00001011110101011110000001100100",
    "10011100100111011011110101111011",
    "00010110001100101001000010100110",
    "11000111000111000000000110011000",
    "11111100100000011110110000111100",
    "10111111111111100101101110100011",
    "11110001101101110100011100101011",
    "01010010000000000011000001000100",
    "01010000110111110001011011001100",
    "00101100111111100111000110010000",
    "11100001111010100111101000111001",
    "01110110101110101001100010110011",
    "10101100011101110101001001010111",
    "01000011000011101111100111001001",
    "10110010100111101011001001001100",
    "00000010001010111101111111111110",
    "11001001001100100110111100001100",
    "01010000111101100111011111111011",
    "11111101110000101000011011101101",
    "00110010011001010000100000100001",
    "10110101110010100001100001001011",
    "11001010111010101110000100010000",
    "00101111110001001011001111100011",
    "01111101000101011010101101101000",
    "00111011010111000001010011111011",
    "00010001101111011110010001110101",
    "01011110100010001011100000010110",
    "01101110111000001111001111000001",
    "11011010011101100000000110111101",
    "00110001100000010101111111110110",
    "10101011000100101001000111011100",
    "11001101001110000001111101110011",
    "00001011011110001010000100110000",
    "11111111101110001110100111111010",
    "00110001111001000010111001010111",
    "00001000110011011101110010111001",
    "11011011111110111000111100001101",
    "00111010001000001100110001110101",
    "00111010100110010001011010011001",
    "00100001000100010100111101110001",
    "10101110010000011000010001001110",
    "10110101001100100101100011110110",
    "00101010100111110010110101100000",
    "00001000010111000101001111110010",
    "11000100111001000001010110001101",
    "01001111001001110010100010110100",
    "00010010000110111001110001001001",
    "01001010100010100100101011101000",
    "11000101100110011111110011111111",
    "00100110100111100100011111011110",
    "00011010011111101001010101001111",
    "01011001001101000100111100111001",
    "00111010101011000010011010011111",
    "00111000101110101111110110101001",
    "01100000011000000110111101000111");

  constant answer_data: output_rom :=(
    "01101101110111110111010011011011",
    "10000000000000000000000000000000",
    "10000000000000000000000000000000",
    "01000111001001001010000100010010",
    "01001000011000100000000011111110",
    "00110101101000000110111100100101",
    "01101010011111001001010000001101",
    "11010011110000111011010011001011",
    "00000111001001101011110100111001",
    "01111001100100010000001011010011",
    "01000111011110111101110001110111",
    "00000001110011100001001001011111",
    "01001001001001010010010101110100",
    "10000000000000000000000000000000",
    "01001010110010011000111001001100",
    "10000000000000000000000000000000",
    "00000000000000000000000000000000",
    "01000101101000101100101000100111",
    "10000001010110101100111001001011",
    "11001000001011101100111011110100",
    "00111001101100011001100010010110",
    "11100011100000000011110110111010",
    "10001001000011110001110101011011",
    "11101011010010110000101011000101",
    "10111101111001101010011010011101",
    "00000000000000000000000000000000",
    "10110100100010000011100010000010",
    "10101100110111101010010110001011",
    "00100001101110011001011111010011",
    "10011001001100110101010001110111",
    "10101011110111100001000100001110",
    "00000000000000000000000000000000",
    "11010111101100010110101010010110",
    "00001110000011100000110101011011",
    "10011001000100101001001111001100",
    "00000000000000000000000000000000",
    "10011000110110001011110011100010",
    "10110111001011101101000001101011",
    "00000000100101001110110000001101",
    "11101100001101001000000100111101",
    "01011101010011001010011101010000",
    "11011000101010000001000001010001",
    "00000000000000000000000000000000",
    "00111100100001000110111110100110",
    "00000000000000000000000000000000",
    "01011110001000101001010111011101",
    "00000000000000000000000000000000",
    "11011111011001100000001110111100",
    "00010001000110011011101001100100",
    "10110000000000100101101100000011",
    "10000000000000000000000000000000",
    "00010101010101100101110101110000",
    "10011010110001101011000011011001",
    "10011111011011011110100001101011",
    "10001000101100010101011110000011",
    "10000000000000000000000000000000",
    "00111001110010011011110101110111",
    "10101111111100010000000110110011",
    "01110010110001000111000100011101",
    "00000000000000000000000000000000",
    "01010111101101001001100011110000",
    "00000100001011110100001111001000",
    "11110110101001011001100000100101",
    "01100110111011011111100011010010",
    "00001110000111001011001001110110",
    "01010010110011011110100101100101",
    "10110110000011000010111001111110",
    "01010010110001110111111101000100",
    "10011011000100011110011010011110",
    "01010011101110010111111110011010",
    "11100000011110010101011100101011",
    "11001111101001011000100100110001",
    "10011101000100000010100010100010",
    "10000000000000000000000000000000",
    "00000100000111100101100110000111",
    "01110010001101100001101000110111",
    "01100011010111110110101011101011",
    "11001111011010010000110101001000",
    "11100011101101000100010101011001",
    "10110110001100010100001101111100",
    "10001011111011111001100010011001",
    "10001111001110110100100011010011",
    "10101000101101001100111000100101",
    "10111011001101000111100101011011",
    "01111001000000001010101110010001",
    "00110000110010101101001111010101",
    "10001001110110000010101111000010",
    "10011101000101000010010011100001",
    "10011001001100101101001001100101",
    "11110010001001001101000111011011",
    "10100101010010100100101001110010",
    "00110101010000000101000011000111",
    "10001111110110111010111111111010",
    "10100000010111011100100110111010",
    "10001101110001000100110101001111",
    "00100001110010110011011101100010",
    "11010000101001100101111011100000",
    "00000001100111010110011110011110",
    "01010100011100101000000011011100",
    "01011001101000111110111100111011");

  signal rom_addr: std_logic_vector(7 downto 0) := (others=>'0');

  signal input1: std_logic_vector(31 downto 0) := (others=>'0');
  signal input2: std_logic_vector(31 downto 0) := (others=>'0');

  signal result1: std_logic_vector(31 downto 0);
  signal result2: std_logic_vector(31 downto 0);

  signal count: std_logic_vector(3 downto 0) := "0000";
  signal errorcount: std_logic_vector(7 downto 0) := "00000000";
  
  signal go : std_logic := '0';
  constant wtime : std_logic_vector(15 downto 0) := x"1B16";--x"362C"; --x"1B16"*2;
  signal writestate : std_logic_vector(3 downto 0) := "1001";
  signal writecountdown : std_logic_vector(15 downto 0) := (others=>'0');
  signal writebuf : std_logic_vector(7 downto 0);

  component fmul
  Port (
    clk    : in  STD_LOGIC;
    input1 : in  STD_LOGIC_VECTOR (31 downto 0);
    input2 : in  STD_LOGIC_VECTOR (31 downto 0);
    output : out STD_LOGIC_VECTOR (31 downto 0));
  end component;

begin
  clk0: clock port map(    
      CLKIN_IN        => MCLK1, 
      RST_IN          => '0', 
      CLKFX_OUT       => clk);

  floatmul: fmul port map(
    clk    => clk,
    input1 => input1,
    input2 => input2,
    output => result1);

  test : process(clk)
  begin
    if rising_edge(clk) then

      result2 <= result1;

      if count < "0011" then
        input1 <= input_data(conv_integer(rom_addr)*2);
        input2 <= input_data(conv_integer(rom_addr)*2 + 1);
        rom_addr <= rom_addr + 1;
        count <= count + 1;

      elsif count = "0011" then
        if rom_addr = 99 then
          count <= "0100";
        end if;
        if answer_data(conv_integer(rom_addr) - 3) /= result2 then
          errorcount <= errorcount + 1;
        end if;
        input1 <= input_data(conv_integer(rom_addr)*2);
        input2 <= input_data(conv_integer(rom_addr)*2 + 1);
        rom_addr <= rom_addr + 1;
        
      elsif count < "0111"  then
        if answer_data(conv_integer(rom_addr) - 3) /= result2 then
          errorcount <= errorcount + 1;
        end if;
        rom_addr <= rom_addr + 1;
        count <= count + 1;
      elsif count = "0111" then
        go <= '1';
        count <= "1111";
      end if;

      if writestate = "1001" then
        if go = '1' then
          RS_TX <= '0';
          writebuf <= errorcount;
          writestate <= "0000";
          writecountdown <= wtime;
        else
          RS_TX <= '1';
        end if;
      elsif writestate = "1000" then
        if writecountdown = 0 then
          RS_TX <= '1';
          writestate <= "1001";
          go <= '0';
        else
          writecountdown <= writecountdown - 1;
        end if;
      else
        if writecountdown = 0 then
          RS_TX <= writebuf(0);
          writebuf <= '1' & writebuf(7 downto 1);
          writecountdown <= wtime;
          writestate <= writestate + 1;
        else
          writecountdown <= writecountdown - 1;
        end if;
      end if;

    end if;
  end process;

end fpu2;

