library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity top is
  Port ( MCLK1 : in  STD_LOGIC;
         RS_TX : out  STD_LOGIC);
end top;

architecture fpu1 of top is

   component clock
    port (
          CLKIN_IN        : in    std_logic; 
          RST_IN          : in    std_logic; 
          CLKFX_OUT       : out   std_logic; 
          CLKIN_IBUFG_OUT : out   std_logic; 
          CLK0_OUT        : out   std_logic; 
          LOCKED_OUT      : out   std_logic);
  end component;

  signal clk: std_logic;
  type input_rom is array(0 to 199) of std_logic_vector(31 downto 0);
  type output_rom is array(0 to 99) of std_logic_vector(31 downto 0);

  constant input_data: input_rom :=(
    "01100111011010010101000101001010",
    "11000110011100111111111111101100",
    "00101001101110101111001011100011",
    "11001101101010111111101101000110",
    "01111100010101000001101111100111",
    "11000010111110001110100010001101",
    "01110110001011100011001111001001",
    "01011010011000111001111110011010",
    "01100110000011010011000110100011",
    "00110010101101110101100001011010",
    "00100101000001010101100001011110",
    "01011101000101111110100111010100",
    "10101011110011011001101101010100",
    "10110010110001101011010000010001",
    "00001110011101000010000111011100",
    "10000010010000010011110110000111",
    "01110000001111100100000111111100",
    "11101001101000011110000101100111",
    "00111110011111101110101001101011",
    "00000001100101111101110010010110",
    "10001111010111001110110000111011",
    "00111000001010101011000011111011",
    "00110010001111001110110011011011",
    "10101111010101000001100001011100",
    "00000010111111101111101110101010",
    "00011010010000111111101000111010",
    "11111011110100010000010101111100",
    "00101001111001100011110010010100",
    "01110101101111101000100101011100",
    "11011000011000011111100110111011",
    "10101000000011111011000111110001",
    "10011001100101011110101110110011",
    "00000101111101111110100100111010",
    "11101111000000001010000111100101",
    "11001010110010110100100001100100",
    "00001011110100000100011110111101",
    "00011111000111100001110001100100",
    "00100011101010000111101111000101",
    "00010100010110100101111001111001",
    "01110011110001010100101101100011",
    "00111011011001000001000100001001",
    "01110000001001001001111011011100",
    "10101010101011000001101110101111",
    "11010100111100100001000000111011",
    "00110011111000110100100000010101",
    "11001101010100000100011101011100",
    "10111011001000101011101001111101",
    "01101111000110011001101111110101",
    "00001011000110100111111111111000",
    "11100001000111000010001100101001",
    "11111000000110111011010101001110",
    "10100100000100111100101011101000",
    "10011000001110000111100100111101",
    "00110010111000000100110100110100",
    "10111100010011101111101001101100",
    "01011111011101111100101100000101",
    "10101100001000011010101001010101",
    "10000110001010110001101010100010",
    "10111110101101010011101101011100",
    "01110000011100110000010011010011",
    "00110110101100111110001011100100",
    "10010100101011111111000010011110",
    "01001111000101011111110101001110",
    "00110010010010011000001010101001",
    "00001000110101001000101001010100",
    "01110000101100100010100101001000",
    "10011010101111000000111010101000",
    "00001010110101010001100001000100",
    "10101100111100110100110000101101",
    "01011011100011101101011110011011",
    "00001001111001011100010010101111",
    "01000010000001100011001111001101",
    "10100011011111111010110101110110",
    "10000100001011011101010001000111",
    "11011110000111000100101000110000",
    "00110010111011001100010011110110",
    "00100000100001011111101100000111",
    "00100011011011001011001000000100",
    "11110100000010110010000010000110",
    "11101100101110011011101011000011",
    "00111110111100011101100100110011",
    "00000101111011000110011110110111",
    "10011001101000110001010011011001",
    "01010000111000111101001100110100",
    "11110111101000000001000011110110",
    "01011110111100101010100000000101",
    "10010100101111101011110001111000",
    "00000001101101000100010011111010",
    "01001001111001101101000011011010",
    "01101001001000110001101001101001",
    "01101010010011000101000110110011",
    "01111110011111100010010101001000",
    "10000100001110101111101110011001",
    "01010011100101000011000110010000",
    "00110010010001001001101111101001",
    "01010111111011101011110011100101",
    "00100101000010001110100101011110",
    "11001111111101011110001001010011",
    "01100000110100101101000011111010",
    "10101010101100101000010101010100",
    "11011000111010000110011001100100",
    "00110101110101001000001010011000",
    "11011001100001110110010101011010",
    "10101000011101010111000010001010",
    "00111111100000000100010001111100",
    "01100010001010011101111010100101",
    "10001001010101111101001110101101",
    "01001110010110010101000110101100",
    "10000110100000000001011110000101",
    "10010101111011001110010011110001",
    "10001100011001100111110001111100",
    "00001100111100011100000010111011",
    "00100010111001001101101000001011",
    "11111100011001100110000101100011",
    "10101111101111001011010000101111",
    "01100010100000110110100100111010",
    "11111111001001111001001100000111",
    "10101111000101101010110000011111",
    "10111000000100010010110111101111",
    "01101101001101001000110101001111",
    "10001001101101100011010111000111",
    "11010100011000111100000111100100",
    "00100100011001111110110100010010",
    "10000011110110001001011011101100",
    "01000101000000101110010111111000",
    "00111001110110000000101010011101",
    "01110111110100011001011011110100",
    "00001001101001011100000100011111",
    "10010101100000100110110010101110",
    "10101010110010100100100110010000",
    "11001101011010001010110010100110",
    "00010110101110100111101011110010",
    "10110100110010101011001000110111",
    "10101000100110011100001000101010",
    "11001011110011111100100110000000",
    "00001000011000011100001101011110",
    "01101110001010000100110001101010",
    "00000011110110101101011100011001",
    "11101101110100110100110010001011",
    "11010010100110010111100100000000",
    "00100010100110100001100011111110",
    "01010110110101001101000111100100",
    "11011001010001011001000100000001",
    "11001101101000111100011011111111",
    "11001001110110010000000100101111",
    "00101010000101010100001111101110",
    "00010101100001110111110001100010",
    "00000010011000010001001110011110",
    "01101001011100101100110101100101",
    "11111100100000010111000110100110",
    "00111110010010010111000111001110",
    "10101011110011110100101100111010",
    "01110101010011111110101001100100",
    "10100111011101100111111011111111",
    "10000001011000011111111010011011",
    "11101011111111011100001101100111",
    "10111111111010010111111000110010",
    "00001101100011000100111010111101",
    "11111001100011001100011110100100",
    "01111100011010100101101100111100",
    "00000010101100100111001011101100",
    "11110100111011010001011011110011",
    "00000001111100000001000001100111",
    "01001101000000001000101111001111",
    "10011001010110111001111111010100",
    "01010000000101111000111010011000",
    "00001010000000111011110000001101",
    "01100001110100011010011110111110",
    "10011011101010111101010100000001",
    "10111111000011101001100011010110",
    "11100101110101100111110111000101",
    "11110010111101100011111000010110",
    "10001110001011101010111111000110",
    "00100001001011010000001010111001",
    "01100011100010100111000011011110",
    "11001001000111111001011100001100",
    "01010110000110100010000100000001",
    "10001001001010110001101100000111",
    "00001101111111010001011010100001",
    "11011000100010111100001010100100",
    "11100011110100101101001001001011",
    "11001111100100101001100000110101",
    "01100001010101010110110011011101",
    "11010101110100010011001111000010",
    "10111100111011010001001111100101",
    "11110111110111101110111100100000",
    "11000111101010111010010010000001",
    "11100010110111010100110110001000",
    "00011100000110101110101100100100",
    "01010011111011100110011001001100",
    "00111011000111101010110001101010",
    "01111001101010001111101101101000",
    "11110011010001100100011100100110",
    "01011000000001100010101100001110",
    "00001101111010110001111100111010",
    "11010010101100100110110000111011",
    "11000000001010101011101011111000",
    "01010100101010110100111011110110",
    "11000111100111100001000111011011",
    "00010110011100110000100000000100");

  constant answer_data: output_rom :=(
    "01100111011010010101000101001010",
    "11001101101010111111101101000110",
    "01111100010101000001101111100111",
    "01110110001011100011001111001001",
    "01100110000011010011000110100011",
    "01011101000101111110100111010100",
    "10110010110001101011011101000111",
    "00001110011101000010000111011100",
    "01110000001111100011110011101101",
    "00111110011111101110101001101011",
    "00111000001010101011000011111011",
    "00110010001110011001110001111010",
    "00011010010000111111101000111010",
    "11111011110100010000010101111100",
    "01110101101111101000100101011100",
    "10101000000011111011000111110001",
    "11101111000000001010000111100101",
    "11001010110010110100100001100100",
    "00100011101010001100101011010011",
    "01110011110001010100101101100011",
    "01110000001001001001111011011100",
    "11010100111100100001000000111011",
    "11001101010100000100011101011100",
    "01101111000110011001101111110101",
    "11100001000111000010001100101001",
    "11111000000110111011010101001110",
    "00110010111000000100110100110100",
    "01011111011101111100101100000101",
    "10101100001000011010101001010101",
    "01110000011100110000010011010011",
    "00110110101100111110001011100100",
    "01001111000101011111110101001110",
    "01110000101100100010100101001000",
    "10011010101111000000111010101000",
    "01011011100011101101011110011011",
    "01000010000001100011001111001101",
    "10100011011111111010110101110110",
    "11011110000111000100101000110000",
    "00100011011100001110000111011100",
    "11110100000010110010000111111001",
    "00111110111100011101100100110011",
    "01010000111000111101001100110100",
    "11110111101000000001000011110110",
    "10010100101111101011110001111000",
    "01101001001000110001101001101001",
    "01111110011111100010010101001000",
    "01010011100101000011000110010000",
    "01010111111011101011110011100101",
    "11001111111101011110001001010011",
    "01100000110100101101000011111010",
    "11011000111010000110011001100100",
    "11011001100001110110010101011010",
    "01100010001010011101111010100101",
    "01001110010110010101000110101100",
    "10010101111011001110010011110001",
    "00001100011111010000010011111010",
    "11111100011001100110000101100011",
    "01100010100000110110100100111010",
    "11111111001001111001001100000111",
    "01101101001101001000110101001111",
    "11010100011000111100000111100100",
    "00100100011001111110110100010010",
    "01000101000000101110010111111001",
    "01110111110100011001011011110100",
    "10101010110010100100100110010000",
    "11001101011010001010110010100110",
    "10110100110010101011001000110111",
    "11001011110011111100100110000000",
    "01101110001010000100110001101010",
    "11101101110100110100110010001011",
    "01010110110101001101000111100100",
    "11011001010001011001000100000010",
    "11001001110110010000000100101111",
    "00010101100001110111110001100010",
    "11111100100000010111000110100110",
    "00111110010010010111000111001110",
    "01110101010011111110101001100100",
    "11101011111111011100001101100111",
    "10111111111010010111111000110010",
    "01111100011001011111010011111111",
    "11110100111011010001011011110011",
    "01001101000000001000101111001111",
    "01010000000101111000111010011000",
    "01100001110100011010011110111110",
    "10111111000011101001100011010110",
    "11110010111101100011111000010110",
    "00100001001011010000001010111001",
    "01100011100010100111000011011110",
    "01010110000110100010000100000001",
    "11011000100010111100001010100100",
    "11100011110100101101001001001011",
    "01100001010101010110110011011100",
    "11110111110111101110111100100000",
    "11100010110111010100110110001000",
    "01010011111011100110011001001100",
    "01111001101010001111101101101000",
    "11110011010001100100011100100110",
    "11010010101100100110110000111011",
    "01010100101010110100111011110110",
    "11000111100111100001000111011011");

  signal rom_addr: std_logic_vector(7 downto 0) := (others=>'0');

  signal input1: std_logic_vector(31 downto 0) := (others=>'0');
  signal input2: std_logic_vector(31 downto 0) := (others=>'0');

  signal result1: std_logic_vector(31 downto 0);
  signal result2: std_logic_vector(31 downto 0);

  signal count: std_logic_vector(3 downto 0) := "0000";
  signal errorcount: std_logic_vector(7 downto 0) := "00000000";
  
  signal go : std_logic := '0';
  constant wtime : std_logic_vector(15 downto 0) := x"362C";
  signal writestate : std_logic_vector(3 downto 0) := "1001";
  signal writecountdown : std_logic_vector(15 downto 0) := (others=>'0');
  signal writebuf : std_logic_vector(7 downto 0);

  component fadd
  Port (
    clk    : in  STD_LOGIC;
    input1 : in  STD_LOGIC_VECTOR (31 downto 0);
    input2 : in  STD_LOGIC_VECTOR (31 downto 0);
    output : out STD_LOGIC_VECTOR (31 downto 0));
  end component;

begin
  clk0: clock port map(    
      CLKIN_IN        => MCLK1, 
      RST_IN          => '0', 
      CLKFX_OUT       => clk);

  floatadd: fadd port map(
    clk    => clk,
    input1 => input1,
    input2 => input2,
    output => result1);

  test : process(clk)
  begin
    if rising_edge(clk) then

      result2 <= result1;

      if count < "0011" then
        input1 <= input_data(conv_integer(rom_addr)*2);
        input2 <= input_data(conv_integer(rom_addr)*2 + 1);
        rom_addr <= rom_addr + 1;
        count <= count + 1;

      elsif count = "0011" then
        if rom_addr = 99 then
          count <= "0100";
        end if;
        if answer_data(conv_integer(rom_addr) - 3) /= result2 then
          errorcount <= errorcount + 1;
        end if;
        input1 <= input_data(conv_integer(rom_addr)*2);
        input2 <= input_data(conv_integer(rom_addr)*2 + 1);
        rom_addr <= rom_addr + 1;
        
      elsif count < "0111"  then
        if answer_data(conv_integer(rom_addr) - 3) /= result2 then
          errorcount <= errorcount + 1;
        end if;
        rom_addr <= rom_addr + 1;
        count <= count + 1;
      elsif count = "0111" then
        go <= '1';
        count <= "1111";
      end if;

      if writestate = "1001" then
        if go = '1' then
          RS_TX <= '0';
          writebuf <= errorcount;
          writestate <= "0000";
          writecountdown <= wtime;
        else
          RS_TX <= '1';
        end if;
      elsif writestate = "1000" then
        if writecountdown = 0 then
          RS_TX <= '1';
          writestate <= "1001";
          go <= '0';
        else
          writecountdown <= writecountdown - 1;
        end if;
      else
        if writecountdown = 0 then
          RS_TX <= writebuf(0);
          writebuf <= '1' & writebuf(7 downto 1);
          writecountdown <= wtime;
          writestate <= writestate + 1;
        else
          writecountdown <= writecountdown - 1;
        end if;
      end if;

    end if;
  end process;

end fpu1;

