library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity top is
  Port ( MCLK1 : in  STD_LOGIC;
         RS_TX : out  STD_LOGIC);
end top;

architecture fpu5 of top is

   component clock
    port (
          CLKIN_IN        : in    std_logic; 
          RST_IN          : in    std_logic; 
          CLKFX_OUT       : out   std_logic; 
          CLKIN_IBUFG_OUT : out   std_logic; 
          CLK0_OUT        : out   std_logic; 
          LOCKED_OUT      : out   std_logic);
  end component;

  signal clk: std_logic;
  type input_rom  is array(0 to 99) of std_logic_vector(31 downto 0);
  type output_rom is array(0 to 99) of std_logic_vector(31 downto 0);

  constant input_data: input_rom :=(
    "01100111110001100110100101110011",
    "01010001111111110100101011101100",
    "00101001110011011011101010101011",
    "11110010111110111110001101000110",
    "01111100110000100101010011111000",
    "00011011111010001110011110001101",
    "01110110010110100010111001100011",
    "00110011100111111100100110011010",
    "01100110001100100000110110110111",
    "00110001010110001010001101011010",
    "00100101010111010000010100010111",
    "01011000111010010101111011010100",
    "10101011101100101100110111000110",
    "10011011101101000101010000010001",
    "00001110100000100111010001000001",
    "00100001001111011101110010000111",
    "01110000111010010011111010100001",
    "01000001111000011111110001100111",
    "00111110000000010111111010010111",
    "11101010110111000110101110010110",
    "10001111001110000101110000101010",
    "11101100101100000011101111111011",
    "00110010101011110011110001010100",
    "11101100000110001101101101011100",
    "00000010000110101111111001000011",
    "11111011111110101010101000111010",
    "11111011001010011101000111100110",
    "00000101001111000111110010010100",
    "01110101110110001011111001100001",
    "10001001111110010101110010111011",
    "10101000100110010000111110010101",
    "10110001111010111111000110110011",
    "00000101111011111111011100000000",
    "11101001101000010011101011100101",
    "11001010000010111100101111010000",
    "01001000010001110110010010111101",
    "00011111001000110001111010101000",
    "00011100011110110110010011000101",
    "00010100011100110101101011000101",
    "01011110010010110111100101100011",
    "00111011011100000110010000100100",
    "00010001100111100000100111011100",
    "10101010110101001010110011110010",
    "00011011000100001010111100111011",
    "00110011110011011110001101010000",
    "01001000010001110001010101011100",
    "10111011011011110010001000011001",
    "10111010100110110111110111110101",
    "00001011111000010001101000011100",
    "01111111001000111111100000101001",
    "11111000101001000001101100010011",
    "10110101110010100100111011101000",
    "10011000001100100011100011100000",
    "01111001010011010011110100110100",
    "10111100010111110100111001110111",
    "11111010110010110110110000000101",
    "10101100100001100010000100101011",
    "10101010000110100101010110100010",
    "10111110011100001011010101110011",
    "00111011000001000101110011010011",
    "00110110100101001011001110101111",
    "11100010111100001110010010011110",
    "01001111001100100001010101001001",
    "11111101100000100100111010101001",
    "00001000011100001101010010110010",
    "10001010001010010101010001001000",
    "10011010000010101011110011010101",
    "00001110000110001010100001000100",
    "10101100010110111111001110001110",
    "01001100110101110010110110011011",
    "00001001010000101110010100000110",
    "11000100001100111010111111001101",
    "10100011100001000111111100101101",
    "10101101110101000111011001000111",
    "11011110001100100001110011101100",
    "01001010110001000011000011110110",
    "00100000001000111000010101101100",
    "11111011101100100000011100000100",
    "11110100111011000000101110111001",
    "00100000101110101000011011000011",
    "00111110000001011111000111101100",
    "11011001011001110011001110110111",
    "10011001010100001010001111100011",
    "00010100110100111101100100110100",
    "11110111010111101010000011110010",
    "00010000101010001111011000000101",
    "10010100000000011011111010110100",
    "10111100010001000111100011111010",
    "01001001011010011110011000100011",
    "11010000000110101101101001101001",
    "01101010011111100100110001111110",
    "01010001001001011011001101001000",
    "10000100010100110011101010010100",
    "11111011001100011001100110010000",
    "00110010010101110100010011101110",
    "10011011101111001110100111100101",
    "00100101110011110000100011110101",
    "11101001111000100101111001010011",
    "01100000101010101101001010110010",
    "11010000100001011111101001010100");

  constant answer_data: output_rom :=(
    "01001110110011111000110011010011",
    "01001110101000111111111010010110",
    "01001110001001110011011011101011",
    "11001101010100000100000111001100",
    "01001110111110011000010010101010",
    "01001101110111110100011100111100",
    "01001110111011001011010001011101",
    "01001110010011100111111100100110",
    "01001110110011000110010000011011",
    "01001110010001010110001010001101",
    "01001110000101010111010000010100",
    "01001110101100011101001010111110",
    "11001110101010001001101001100100",
    "11001110110010001001011101011000",
    "01001101011010000010011101000100",
    "01001110000001001111011101110010",
    "01001110111000011101001001111101",
    "01001110100000111100001111111001",
    "01001110011110000000010111111010",
    "11001101101010010001110010100011",
    "11001110111000011000111101001000",
    "11001101100110100111111000100000",
    "01001110010010101011110011110001",
    "11001101100111110011100100100101",
    "01001100000001101011111110010001",
    "11001100100000001010101010111001",
    "11001100100110101100010111000011",
    "01001100101001111000111110010011",
    "01001110111010111011000101111101",
    "11001110111011000000110101000111",
    "11001110101011101100110111100001",
    "11001110100111000010100000011101",
    "01001100101111011111111011100000",
    "11001101101100101111011000101001",
    "11001110010101111101000011010001",
    "01001110100100001000111011001001",
    "01001101111110010001100011110101",
    "01001101111000111101101100100110",
    "01001101101000111001101011010110",
    "01001110101111001001011011110011",
    "01001110011011011100000110010001",
    "01001101100011001111000001001111",
    "11001110101010100101011010100110",
    "01001101110110001000010101111010",
    "01001110010011110011011110001101",
    "01001110100100001000111000101011",
    "11001110100010010010000110111100",
    "11001110100010101100100100000100",
    "01001101001111100001000110100010",
    "01001110111111100100011111110000",
    "11001100111010110111110010011110",
    "11001110100101000110101101100010",
    "11001110110011111001101110001110",
    "01001110111100101001101001111010",
    "11001110100001110100000101100011",
    "11001100101001101001001001111111",
    "11001110101001101111001110111110",
    "11001110101010111100101101010101",
    "11001110100000110001111010010101",
    "01001110011011000001000101110011",
    "01001110010110100101001011001111",
    "11001101111010000111100011011011",
    "01001110100111100110010000101011",
    "11001100000111110110110001010110",
    "01001101000001110000110101001011",
    "11001110111010111010110101010111",
    "11001110110010111110101010000110",
    "01001101011000011000101010000100",
    "11001110101001110100100000011001",
    "01001110100110011010111001011011",
    "01001101000101000010111001010000",
    "11001110011011110011000101000001",
    "11001110101110001111011100000010",
    "11001110101001000101011100010011",
    "11001110000001110011011110001100",
    "01001110100101011000100001100010",
    "01001110000000001000111000010110",
    "11001100100010011011111100100000",
    "11001101001100010011111101000100",
    "01001110000000101110101000011011",
    "01001110011110000001011111001000",
    "11001110000110100110001100110001",
    "11001110110011010101111010111000",
    "01001101101001101001111011001010",
    "11001101000010100001010111110001",
    "01001101100001010100011110110000",
    "11001110110101111111110010000011",
    "11001110100001110111011100001110",
    "01001110100100101101001111001100",
    "11001110001111111001010010010110",
    "01001110110101001111110010011001",
    "01001110101000100100101101100111",
    "11001110111101110101100110001011",
    "11001100100110011100110011001110",
    "01001110010010010101110100010100",
    "11001110110010001000011000101100",
    "01001110000101110011110000100100",
    "11001101101100001110110100001101",
    "01001110110000010101010110100101",
    "11001110001111011110100000010111");

  signal rom_addr: std_logic_vector(7 downto 0) := (others=>'0');
  signal input: std_logic_vector(31 downto 0) := (others=>'0');
  signal result1: std_logic_vector(31 downto 0);
  signal result2: std_logic_vector(31 downto 0);
  signal count: std_logic_vector(3 downto 0) := "0000";
  signal errorcount: std_logic_vector(7 downto 0) := "00000000";
  signal go : std_logic := '0';
  constant wtime : std_logic_vector(15 downto 0) := x"362C";
  signal writestate : std_logic_vector(3 downto 0) := "1001";
  signal writecountdown : std_logic_vector(15 downto 0) := (others=>'0');
  signal writebuf : std_logic_vector(7 downto 0);

  component itof
  Port (
    clk    : in  STD_LOGIC;
    input  : in  STD_LOGIC_VECTOR (31 downto 0);
    output : out STD_LOGIC_VECTOR (31 downto 0));
  end component;

begin
  clk0: clock port map(    
      CLKIN_IN        => MCLK1, 
      RST_IN          => '0', 
      CLKFX_OUT       => clk);

  inttofloat: itof port map(
    clk    => clk,
    input  => input,
    output => result1);

  test : process(clk)
  begin
    if rising_edge(clk) then

      result2 <= result1;

      if count < "0011" then
        input <= input_data(conv_integer(rom_addr));
        rom_addr <= rom_addr + 1;
        count <= count + 1;

      elsif count = "0011" then
        if rom_addr = 99 then
          count <= "0100";
        end if;
        if answer_data(conv_integer(rom_addr) - 3) /= result2 then
          errorcount <= errorcount + 1;
        end if;
        input <= input_data(conv_integer(rom_addr));
        rom_addr <= rom_addr + 1;
        
      elsif count < "0111"  then
        if answer_data(conv_integer(rom_addr) - 3) /= result2 then
          errorcount <= errorcount + 1;
        end if;
        rom_addr <= rom_addr + 1;
        count <= count + 1;
      elsif count = "0111" then
        go <= '1';
        count <= "1111";
      end if;


      if writestate = "1001" then
        if go = '1' then
          RS_TX <= '0';
          writebuf <= errorcount;
          writestate <= "0000";
          writecountdown <= wtime;
        else
          RS_TX <= '1';
        end if;
      elsif writestate = "1000" then
        if writecountdown = 0 then
          RS_TX <= '1';
          writestate <= "1001";
          go <= '0';
        else
          writecountdown <= writecountdown - 1;
        end if;
      else
        if writecountdown = 0 then
          RS_TX <= writebuf(0);
          writebuf <= '1' & writebuf(7 downto 1);
          writecountdown <= wtime;
          writestate <= writestate + 1;
        else
          writecountdown <= writecountdown - 1;
        end if;
      end if;

    end if;
  end process;

end fpu5;

