-- TestBench Template

  LIBRARY ieee;
  USE ieee.std_logic_1164.ALL;
  USE ieee.numeric_std.ALL;

  use work.types.all;

  ENTITY testbench IS
      generic (
          wtime : std_logic_vector (15 downto 0) := x"0010"
      );
  END testbench;

  ARCHITECTURE behavior OF testbench IS

  -- Component Declaration
          COMPONENT TOP
          generic (
--              wtime : std_logic_vector (15 downto 0) := x"1ADB"
              wtime : std_logic_vector (15 downto 0) := wtime
          );
          PORT(
                  MCLK1 : in std_logic;
                  RS_RX : in std_logic;
                  RS_TX : out std_logic;
                  ZD     : inout std_logic_vector (31 downto 0);
                  ZA     : out   std_logic_vector (19 downto 0);
                  XWA    : out   std_logic;
                  XE1    : out   std_logic;
                  E2A    : out   std_logic;
                  XE3    : out   std_logic;
                  XGA    : out   std_logic;
                  XZCKE  : out   std_logic;
                  ADVA   : out   std_logic;
                  XLBO   : out   std_logic;
                  ZZA    : out   std_logic;
                  XFT    : out   std_logic;
                  XZBE   : out   std_logic_vector (3 downto 0);
                  ZCLKMA : out   std_logic_vector (1 downto 0));
          END COMPONENT;
          component sram_sim port (
                  ZD     : inout std_logic_vector (31 downto 0);
                  ZA     : in std_logic_vector (19 downto 0);
                  XWA    : in std_logic;
                  XE1    : in std_logic;
                  E2A    : in std_logic;
                  XE3    : in std_logic;
                  XGA    : in std_logic;
                  XZCKE  : in std_logic;
                  ADVA   : in std_logic;
                  XLBO   : in std_logic;
                  ZZA    : in std_logic;
                  XFT    : in std_logic;
                  XZBE   : in std_logic_vector (3 downto 0);
                  ZCLKMA : in std_logic_vector (1 downto 0));
          end component;
          signal clk : std_logic;
          signal rs_rx : std_logic;
          signal rs_tx : std_logic;
          signal zd     : std_logic_vector (31 downto 0);
          signal za     : std_logic_vector (19 downto 0);
          signal xwa    : std_logic;
          signal xe1    : std_logic;
          signal e2a    : std_logic;
          signal xe3    : std_logic;
          signal xga    : std_logic;
          signal xzcke  : std_logic;
          signal adva   : std_logic;
          signal xlbo   : std_logic;
          signal zza    : std_logic;
          signal xft    : std_logic;
          signal xzbe   : std_logic_vector (3 downto 0);
          signal zclkma : std_logic_vector (1 downto 0);
          signal rst : std_logic := '0';
          signal receiver_in : receiver_in_type;
          signal receiver_out : receiver_out_type;
          signal sender_in : sender_in_type;
          signal sender_out : sender_out_type;
          signal counter : std_logic_vector (15 downto 0) := x"b284";
          type inst_list_type is array (45700 downto 0) of std_logic_vector (7 downto 0);
          signal inst_list : inst_list_type := (
x"02", x"00", x"00", x"39", 
x"40", x"c9", x"0f", x"db", 
x"40", x"49", x"0f", x"db", 
x"3f", x"c9", x"0f", x"db", 
x"3f", x"49", x"0f", x"db", 
x"3f", x"80", x"00", x"00", 
x"40", x"00", x"00", x"00", 
x"bf", x"80", x"00", x"00", 
x"3f", x"00", x"00", x"00", 
x"3d", x"cc", x"cc", x"cd", 
x"cb", x"00", x"00", x"00", 
x"4b", x"00", x"00", x"00", 
x"bf", x"00", x"00", x"00", 
x"3d", x"2a", x"a7", x"89", 
x"ba", x"b3", x"81", x"06", 
x"be", x"2a", x"aa", x"ac", 
x"3c", x"08", x"86", x"66", 
x"b9", x"4d", x"64", x"b6", 
x"3e", x"e0", x"00", x"00", 
x"40", x"1c", x"00", x"00", 
x"be", x"aa", x"aa", x"aa", 
x"3e", x"4c", x"cc", x"cd", 
x"be", x"12", x"49", x"25", 
x"3d", x"e3", x"8e", x"38", 
x"bd", x"b7", x"d6", x"6e", 
x"3d", x"75", x"e7", x"c5", 
x"43", x"00", x"00", x"00", 
x"3f", x"66", x"66", x"66", 
x"3e", x"4c", x"cc", x"cd", 
x"43", x"16", x"00", x"00", 
x"c3", x"16", x"00", x"00", 
x"3d", x"cc", x"cc", x"cd", 
x"c0", x"00", x"00", x"00", 
x"3b", x"80", x"00", x"00", 
x"41", x"a0", x"00", x"00", 
x"3d", x"4c", x"cc", x"cd", 
x"3e", x"80", x"00", x"00", 
x"41", x"20", x"00", x"00", 
x"3e", x"99", x"99", x"9a", 
x"43", x"7f", x"00", x"00", 
x"3e", x"19", x"99", x"9a", 
x"40", x"49", x"0f", x"db", 
x"41", x"f0", x"00", x"00", 
x"41", x"70", x"00", x"00", 
x"38", x"d1", x"b7", x"17", 
x"4c", x"be", x"bc", x"20", 
x"4e", x"6e", x"6b", x"28", 
x"bd", x"cc", x"cc", x"cd", 
x"3c", x"23", x"d7", x"0a", 
x"be", x"4c", x"cc", x"cd", 
x"3f", x"00", x"00", x"00", 
x"40", x"00", x"00", x"00", 
x"c3", x"48", x"00", x"00", 
x"43", x"48", x"00", x"00", 
x"3c", x"8e", x"fa", x"35", 
x"bf", x"80", x"00", x"00", 
x"3f", x"80", x"00", x"00", 
x"00", x"00", x"00", x"00", 
x"01", x"00", x"2c", x"65", 
x"08", x"20", x"00", x"aa", 
x"74", x"20", x"00", x"00", 
x"20", x"00", x"26", x"33", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"18", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"18", x"00", 
x"84", x"42", x"18", x"00", 
x"94", x"42", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"64", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"80", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"20", x"80", x"00", x"18", 
x"08", x"60", x"00", x"37", 
x"c0", x"43", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"20", x"60", x"00", x"1a", 
x"08", x"60", x"00", x"36", 
x"c0", x"63", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"63", x"10", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a5", x"10", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"84", x"a5", x"10", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"20", x"00", 
x"84", x"45", x"10", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"62", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"82", x"20", x"00", 
x"84", x"63", x"20", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"08", x"a0", x"00", x"01", 
x"07", x"62", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"82", x"20", x"00", 
x"84", x"63", x"20", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"08", x"a0", x"00", x"02", 
x"07", x"62", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"42", x"20", x"00", 
x"84", x"63", x"10", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"62", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"08", x"a0", x"00", x"01", 
x"07", x"62", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"08", x"a0", x"00", x"02", 
x"07", x"62", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"62", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"08", x"c0", x"00", x"01", 
x"07", x"62", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"08", x"c0", x"00", x"02", 
x"07", x"62", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"c0", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"50", x"00", x"05", 
x"40", x"70", x"00", x"04", 
x"40", x"90", x"00", x"03", 
x"40", x"b0", x"00", x"02", 
x"40", x"d0", x"00", x"01", 
x"08", x"e0", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"a4", x"ff", x"fe", 
x"47", x"a5", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"a7", x"ff", x"fb", 
x"47", x"a6", x"ff", x"fa", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"47", x"a2", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"5d", x"ff", x"f9", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"47", x"a2", x"ff", x"f8", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"c7", x"a2", x"ff", x"f7", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"c0", x"7d", x"ff", x"f7", 
x"c7", x"a2", x"ff", x"f6", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"c7", x"a2", x"ff", x"f5", 
x"0b", x"bd", x"ff", x"f4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0c", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"c7", x"a2", x"ff", x"f4", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"c0", x"7d", x"ff", x"f4", 
x"c7", x"a2", x"ff", x"f3", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"c0", x"7d", x"ff", x"f6", 
x"8c", x"83", x"10", x"00", 
x"08", x"60", x"00", x"34", 
x"c0", x"a3", x"00", x"00", 
x"8c", x"84", x"28", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"80", x"00", x"33", 
x"c0", x"84", x"00", x"00", 
x"c0", x"bd", x"ff", x"f5", 
x"8c", x"85", x"20", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"c0", x"9d", x"ff", x"f3", 
x"8c", x"c3", x"20", x"00", 
x"08", x"80", x"00", x"34", 
x"c0", x"e4", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"a0", x"00", x"38", 
x"c0", x"c5", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"98", x"c2", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"98", x"c5", x"00", x"00", 
x"8c", x"c6", x"10", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"10", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"98", x"63", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"98", x"a5", x"00", x"00", 
x"8c", x"a5", x"20", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"07", x"65", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"40", x"9d", x"ff", x"ff", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"50", x"00", x"02", 
x"40", x"70", x"00", x"01", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"c7", x"a2", x"ff", x"fd", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"40", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"c0", x"7d", x"ff", x"fd", 
x"c7", x"a2", x"ff", x"fc", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"c0", x"7d", x"ff", x"fc", 
x"c7", x"a2", x"ff", x"fb", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"00", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"43", x"10", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"c0", x"5d", x"ff", x"fc", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"02", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"47", x"a2", x"ff", x"fa", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c7", x"a2", x"ff", x"fd", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c7", x"a2", x"ff", x"fc", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c7", x"a2", x"ff", x"fb", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c7", x"a2", x"ff", x"fa", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c7", x"a2", x"ff", x"f9", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"c0", x"7d", x"ff", x"f9", 
x"c0", x"9d", x"ff", x"fb", 
x"8c", x"a4", x"18", x"00", 
x"c0", x"dd", x"ff", x"fa", 
x"c0", x"fd", x"ff", x"fc", 
x"8d", x"07", x"30", x"00", 
x"8d", x"08", x"18", x"00", 
x"c1", x"3d", x"ff", x"fd", 
x"8d", x"49", x"10", x"00", 
x"89", x"08", x"50", x"00", 
x"8d", x"49", x"30", x"00", 
x"8d", x"4a", x"18", x"00", 
x"8d", x"67", x"10", x"00", 
x"85", x"4a", x"58", x"00", 
x"8d", x"64", x"10", x"00", 
x"8d", x"87", x"30", x"00", 
x"8d", x"8c", x"10", x"00", 
x"8d", x"a9", x"18", x"00", 
x"85", x"8c", x"68", x"00", 
x"8d", x"a9", x"30", x"00", 
x"8d", x"ad", x"10", x"00", 
x"8c", x"67", x"18", x"00", 
x"89", x"ad", x"18", x"00", 
x"98", x"c6", x"00", x"00", 
x"8c", x"e7", x"20", x"00", 
x"8d", x"29", x"20", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"63", x"10", x"00", 
x"c0", x"9b", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"8d", x"c5", x"28", x"00", 
x"8d", x"c2", x"70", x"00", 
x"8d", x"eb", x"58", x"00", 
x"8d", x"e3", x"78", x"00", 
x"85", x"ce", x"78", x"00", 
x"8d", x"e6", x"30", x"00", 
x"8d", x"e4", x"78", x"00", 
x"85", x"ce", x"78", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"6e", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"8d", x"c8", x"40", x"00", 
x"8d", x"c2", x"70", x"00", 
x"8d", x"ec", x"60", x"00", 
x"8d", x"e3", x"78", x"00", 
x"85", x"ce", x"78", x"00", 
x"8d", x"e7", x"38", x"00", 
x"8d", x"e4", x"78", x"00", 
x"85", x"ce", x"78", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"6e", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"8d", x"ca", x"50", x"00", 
x"8d", x"c2", x"70", x"00", 
x"8d", x"ed", x"68", x"00", 
x"8d", x"e3", x"78", x"00", 
x"85", x"ce", x"78", x"00", 
x"8d", x"e9", x"48", x"00", 
x"8d", x"e4", x"78", x"00", 
x"85", x"ce", x"78", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"6e", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"32", 
x"c1", x"c3", x"00", x"00", 
x"8d", x"e2", x"40", x"00", 
x"8d", x"ef", x"50", x"00", 
x"8e", x"03", x"60", x"00", 
x"8e", x"10", x"68", x"00", 
x"85", x"ef", x"80", x"00", 
x"8e", x"04", x"38", x"00", 
x"8e", x"10", x"48", x"00", 
x"85", x"ef", x"80", x"00", 
x"8d", x"ce", x"78", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c7", x"6e", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"80", x"00", x"32", 
x"c1", x"c4", x"00", x"00", 
x"8d", x"e2", x"28", x"00", 
x"8d", x"ef", x"50", x"00", 
x"8d", x"43", x"58", x"00", 
x"8d", x"4a", x"68", x"00", 
x"85", x"ef", x"50", x"00", 
x"8d", x"44", x"30", x"00", 
x"8d", x"4a", x"48", x"00", 
x"85", x"ef", x"50", x"00", 
x"8d", x"ce", x"78", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"6e", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"80", x"00", x"32", 
x"c1", x"24", x"00", x"00", 
x"8c", x"42", x"28", x"00", 
x"8c", x"42", x"40", x"00", 
x"8c", x"63", x"58", x"00", 
x"8c", x"63", x"60", x"00", 
x"84", x"42", x"18", x"00", 
x"8c", x"84", x"30", x"00", 
x"8c", x"84", x"38", x"00", 
x"84", x"42", x"20", x"00", 
x"8d", x"29", x"10", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"69", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"01", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"5b", x"02", x"52", 
x"47", x"a2", x"ff", x"fd", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"47", x"a2", x"ff", x"fc", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"47", x"a2", x"ff", x"fb", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"47", x"a3", x"ff", x"f9", 
x"47", x"a2", x"ff", x"f8", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"40", x"5d", x"ff", x"f9", 
x"40", x"7d", x"ff", x"f8", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"47", x"a2", x"ff", x"f7", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f8", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"47", x"a2", x"ff", x"f6", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f6", 
x"40", x"7d", x"ff", x"f8", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"60", x"00", x"00", 
x"47", x"a3", x"ff", x"f5", 
x"47", x"a2", x"ff", x"f4", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"40", x"5d", x"ff", x"f5", 
x"40", x"7d", x"ff", x"f4", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"47", x"a2", x"ff", x"f3", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"f4", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"47", x"a2", x"ff", x"f2", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"40", x"5d", x"ff", x"f2", 
x"40", x"7d", x"ff", x"f4", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"f1", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"08", x"60", x"00", x"00", 
x"47", x"a3", x"ff", x"f0", 
x"47", x"a2", x"ff", x"ef", 
x"0b", x"bd", x"ff", x"ee", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"12", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"7d", x"ff", x"ef", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"47", x"a2", x"ff", x"ee", 
x"0b", x"bd", x"ff", x"ed", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"13", 
x"40", x"5d", x"ff", x"ee", 
x"40", x"7d", x"ff", x"ef", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"ed", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"13", 
x"08", x"60", x"00", x"00", 
x"47", x"a3", x"ff", x"ed", 
x"47", x"a2", x"ff", x"ec", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"40", x"5d", x"ff", x"ed", 
x"40", x"7d", x"ff", x"ec", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"47", x"a2", x"ff", x"eb", 
x"0b", x"bd", x"ff", x"ea", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"16", 
x"40", x"5d", x"ff", x"eb", 
x"40", x"7d", x"ff", x"ec", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"47", x"a2", x"ff", x"ea", 
x"0b", x"bd", x"ff", x"e9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"17", 
x"40", x"5d", x"ff", x"ea", 
x"40", x"7d", x"ff", x"ec", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"17", 
x"40", x"7d", x"ff", x"fa", 
x"47", x"a2", x"ff", x"e9", 
x"20", x"60", x"00", x"2b", 
x"08", x"80", x"00", x"00", 
x"47", x"a4", x"ff", x"e8", 
x"0b", x"bd", x"ff", x"e7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"19", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"40", x"5d", x"ff", x"e8", 
x"40", x"7d", x"ff", x"e9", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"47", x"a2", x"ff", x"e7", 
x"0b", x"bd", x"ff", x"e6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1a", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"40", x"5d", x"ff", x"e7", 
x"40", x"7d", x"ff", x"e9", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"47", x"a2", x"ff", x"e6", 
x"0b", x"bd", x"ff", x"e5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"e0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1b", 
x"08", x"40", x"00", x"35", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"40", x"5d", x"ff", x"e6", 
x"40", x"7d", x"ff", x"e9", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"0b", x"60", x"00", x"02", 
x"20", x"5b", x"00", x"02", 
x"40", x"7d", x"ff", x"f1", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"04", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a3", x"ff", x"e5", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"0b", 
x"44", x"62", x"00", x"0a", 
x"40", x"5d", x"ff", x"e9", 
x"44", x"62", x"00", x"09", 
x"40", x"9d", x"ff", x"ec", 
x"44", x"64", x"00", x"08", 
x"40", x"9d", x"ff", x"ef", 
x"44", x"64", x"00", x"07", 
x"40", x"9d", x"ff", x"e5", 
x"44", x"64", x"00", x"06", 
x"40", x"9d", x"ff", x"f4", 
x"44", x"64", x"00", x"05", 
x"40", x"9d", x"ff", x"f8", 
x"44", x"64", x"00", x"04", 
x"40", x"bd", x"ff", x"fa", 
x"44", x"65", x"00", x"03", 
x"40", x"dd", x"ff", x"fb", 
x"44", x"66", x"00", x"02", 
x"40", x"dd", x"ff", x"fc", 
x"44", x"66", x"00", x"01", 
x"40", x"fd", x"ff", x"fd", 
x"44", x"67", x"00", x"00", 
x"40", x"fd", x"ff", x"ff", 
x"41", x"1d", x"ff", x"fe", 
x"07", x"68", x"38", x"00", 
x"47", x"63", x"00", x"00", 
x"0b", x"60", x"00", x"03", 
x"20", x"db", x"00", x"38", 
x"0b", x"60", x"00", x"02", 
x"20", x"db", x"00", x"0c", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"7d", x"ff", x"f1", 
x"20", x"60", x"00", x"14", 
x"08", x"60", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"16", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"40", x"5d", x"ff", x"fa", 
x"20", x"40", x"00", x"09", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"e9", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"16", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"40", x"5d", x"ff", x"fa", 
x"20", x"40", x"00", x"09", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"e9", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"01", 
x"20", x"c0", x"00", x"03", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"20", x"00", x"00", x"17", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"0f", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"ac", x"43", x"00", x"06", 
x"08", x"c0", x"00", x"37", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"20", x"00", x"00", x"05", 
x"08", x"c0", x"00", x"36", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"20", x"00", x"00", x"05", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"01", 
x"20", x"c0", x"00", x"5a", 
x"08", x"c0", x"00", x"38", 
x"c0", x"46", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"3f", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"29", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"ac", x"43", x"00", x"13", 
x"08", x"c0", x"00", x"37", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"36", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"46", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"01", 
x"20", x"c0", x"00", x"03", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"20", x"00", x"00", x"08", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"ac", x"43", x"00", x"03", 
x"08", x"c0", x"00", x"37", 
x"c0", x"66", x"00", x"00", 
x"20", x"00", x"00", x"02", 
x"08", x"c0", x"00", x"36", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"3f", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"a0", x"43", x"00", x"29", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"ac", x"43", x"00", x"13", 
x"08", x"c0", x"00", x"37", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"36", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"10", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"46", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"a0", x"00", x"09", 
x"08", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"02", x"21", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"02", 
x"40", x"90", x"00", x"01", 
x"0b", x"60", x"00", x"3c", 
x"2f", x"62", x"00", x"2f", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"47", x"a4", x"ff", x"fd", 
x"47", x"a2", x"ff", x"fc", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"05", x"3f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"20", x"40", x"00", x"1c", 
x"40", x"5d", x"ff", x"fc", 
x"08", x"42", x"00", x"01", 
x"0b", x"60", x"00", x"3c", 
x"2f", x"62", x"00", x"17", 
x"40", x"7d", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fb", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"05", x"4e", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"20", x"40", x"00", x"06", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"0a", x"03", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"47", x"64", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"47", x"64", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"5b", x"00", x"0e", 
x"40", x"7d", x"ff", x"ff", 
x"08", x"83", x"00", x"01", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"62", x"18", x"00", 
x"47", x"64", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"ff", 
x"08", x"42", x"00", x"01", 
x"08", x"60", x"ff", x"ff", 
x"20", x"00", x"24", x"b0", 
x"08", x"60", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"5b", x"00", x"0e", 
x"40", x"5d", x"ff", x"ff", 
x"08", x"82", x"00", x"01", 
x"47", x"a3", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"7f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"62", x"18", x"00", 
x"47", x"64", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"ff", 
x"08", x"42", x"00", x"01", 
x"20", x"00", x"24", x"91", 
x"40", x"70", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"7b", x"00", x"1b", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"63", x"00", x"01", 
x"08", x"40", x"00", x"00", 
x"47", x"a3", x"ff", x"fc", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"7b", x"00", x"09", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"43", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"0a", x"03", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"50", x"00", x"06", 
x"40", x"70", x"00", x"05", 
x"40", x"90", x"00", x"04", 
x"40", x"b0", x"00", x"03", 
x"40", x"d0", x"00", x"02", 
x"40", x"f0", x"00", x"01", 
x"47", x"a5", x"ff", x"ff", 
x"47", x"a7", x"ff", x"fe", 
x"47", x"a6", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"a4", x"ff", x"fb", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"05", x"db", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"40", x"5d", x"ff", x"fb", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"05", x"e4", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"05", x"ee", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"7b", x"00", x"1c", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"06", x"0a", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"47", x"a2", x"ff", x"f9", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"7f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"7d", x"ff", x"f9", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"47", x"a2", x"ff", x"f9", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"05", x"7f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"7d", x"ff", x"f9", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"f0", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"09", x"00", x"00", x"38", 
x"c0", x"c8", x"00", x"00", 
x"a0", x"a6", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"09", x"00", x"00", x"01", 
x"21", x"00", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"41", x"02", x"00", x"04", 
x"40", x"42", x"00", x"06", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"09", x"20", x"00", x"38", 
x"c0", x"c9", x"00", x"00", 
x"ac", x"c5", x"00", x"02", 
x"09", x"20", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"09", x"20", x"00", x"00", 
x"20", x"40", x"00", x"44", 
x"21", x"20", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"40", x"00", x"01", 
x"07", x"68", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"20", x"40", x"00", x"1e", 
x"88", x"a5", x"10", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"a5", x"d8", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"18", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"0f", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"20", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"67", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"98", x"a5", x"00", x"00", 
x"88", x"a5", x"10", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"a5", x"d8", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"18", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"0f", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"20", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"67", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"07", x"68", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"21", x"20", x"00", x"1e", 
x"88", x"a5", x"10", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"a5", x"d8", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"18", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"0f", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"20", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"67", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"98", x"a5", x"00", x"00", 
x"88", x"a5", x"10", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"a5", x"d8", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"18", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"0f", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"20", x"00", 
x"9c", x"42", x"00", x"00", 
x"07", x"68", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"67", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"08", x"e0", x"00", x"02", 
x"c7", x"a2", x"ff", x"ff", 
x"c7", x"a4", x"ff", x"fe", 
x"c7", x"a3", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"a2", x"ff", x"fb", 
x"47", x"a4", x"ff", x"fa", 
x"0a", x"04", x"00", x"00", 
x"08", x"85", x"00", x"00", 
x"08", x"a6", x"00", x"00", 
x"08", x"c7", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"06", x"d6", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"08", x"a0", x"00", x"02", 
x"08", x"c0", x"00", x"00", 
x"c0", x"5d", x"ff", x"fd", 
x"c0", x"7d", x"ff", x"fe", 
x"c0", x"9d", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"fd", x"ff", x"fa", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"06", x"ea", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"02", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"08", x"a0", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"c0", x"5d", x"ff", x"fe", 
x"c0", x"7d", x"ff", x"ff", 
x"c0", x"9d", x"ff", x"fd", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"fd", x"ff", x"fa", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"06", x"fe", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"03", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"8c", x"a2", x"10", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"8c", x"c3", x"18", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"84", x"a5", x"30", x"00", 
x"8c", x"c4", x"20", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"02", 
x"07", x"63", x"20", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"84", x"a5", x"30", x"00", 
x"40", x"62", x"00", x"03", 
x"20", x"60", x"00", x"16", 
x"8c", x"c3", x"20", x"00", 
x"40", x"62", x"00", x"09", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"84", x"a5", x"30", x"00", 
x"8c", x"84", x"10", x"00", 
x"40", x"62", x"00", x"09", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"84", x"30", x"00", 
x"84", x"a5", x"20", x"00", 
x"8c", x"42", x"18", x"00", 
x"40", x"42", x"00", x"09", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"84", x"45", x"10", x"00", 
x"33", x"e0", x"00", x"00", 
x"80", x"45", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"8d", x"02", x"28", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c1", x"3b", x"00", x"00", 
x"8d", x"08", x"48", x"00", 
x"8d", x"23", x"30", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c1", x"5b", x"00", x"00", 
x"8d", x"29", x"50", x"00", 
x"85", x"08", x"48", x"00", 
x"8d", x"24", x"38", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"02", 
x"07", x"63", x"20", x"00", 
x"c1", x"5b", x"00", x"00", 
x"8d", x"29", x"50", x"00", 
x"85", x"08", x"48", x"00", 
x"40", x"62", x"00", x"03", 
x"20", x"60", x"00", x"1f", 
x"8d", x"24", x"30", x"00", 
x"8d", x"43", x"38", x"00", 
x"85", x"29", x"50", x"00", 
x"40", x"62", x"00", x"09", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c1", x"5b", x"00", x"00", 
x"8d", x"29", x"50", x"00", 
x"8c", x"e2", x"38", x"00", 
x"8c", x"84", x"28", x"00", 
x"84", x"e7", x"20", x"00", 
x"40", x"62", x"00", x"09", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"e7", x"20", x"00", 
x"85", x"29", x"38", x"00", 
x"8c", x"42", x"30", x"00", 
x"8c", x"63", x"28", x"00", 
x"84", x"42", x"18", x"00", 
x"40", x"42", x"00", x"09", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"85", x"29", x"10", x"00", 
x"08", x"40", x"00", x"31", 
x"c0", x"42", x"00", x"00", 
x"8d", x"29", x"10", x"00", 
x"84", x"48", x"48", x"00", 
x"33", x"e0", x"00", x"00", 
x"80", x"48", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"db", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"fb", x"00", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"c7", x"a4", x"ff", x"fe", 
x"c7", x"a3", x"ff", x"fd", 
x"c7", x"a2", x"ff", x"fc", 
x"47", x"a2", x"ff", x"fb", 
x"47", x"a3", x"ff", x"fa", 
x"80", x"87", x"00", x"00", 
x"80", x"66", x"00", x"00", 
x"80", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"05", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"40", x"00", x"01", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"c0", x"9b", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"63", x"10", x"00", 
x"c0", x"bb", x"00", x"00", 
x"c0", x"dd", x"ff", x"fc", 
x"c0", x"fd", x"ff", x"fd", 
x"c1", x"1d", x"ff", x"fe", 
x"40", x"5d", x"ff", x"fb", 
x"c7", x"a2", x"ff", x"f9", 
x"80", x"43", x"00", x"00", 
x"80", x"64", x"00", x"00", 
x"80", x"85", x"00", x"00", 
x"80", x"a6", x"00", x"00", 
x"80", x"c7", x"00", x"00", 
x"80", x"e8", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"33", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"c0", x"7d", x"ff", x"fc", 
x"c0", x"9d", x"ff", x"fd", 
x"c0", x"bd", x"ff", x"fe", 
x"40", x"5d", x"ff", x"fb", 
x"c7", x"a2", x"ff", x"f8", 
x"80", x"43", x"00", x"00", 
x"80", x"64", x"00", x"00", 
x"80", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"05", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"62", x"00", x"01", 
x"0b", x"60", x"00", x"03", 
x"20", x"7b", x"00", x"20", 
x"c0", x"7d", x"ff", x"f8", 
x"8c", x"83", x"18", x"00", 
x"c0", x"bd", x"ff", x"f9", 
x"8c", x"45", x"10", x"00", 
x"88", x"84", x"10", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"ac", x"82", x"00", x"16", 
x"94", x"84", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"09", 
x"08", x"40", x"00", x"00", 
x"88", x"84", x"18", x"00", 
x"93", x"65", x"00", x"00", 
x"8c", x"84", x"d8", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"98", x"84", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"88", x"84", x"18", x"00", 
x"93", x"65", x"00", x"00", 
x"8c", x"84", x"d8", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"c0", x"7d", x"ff", x"f8", 
x"8c", x"83", x"18", x"00", 
x"c0", x"bd", x"ff", x"f9", 
x"8c", x"45", x"10", x"00", 
x"88", x"84", x"10", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"ac", x"82", x"00", x"16", 
x"94", x"84", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"09", 
x"08", x"40", x"00", x"00", 
x"88", x"84", x"18", x"00", 
x"93", x"65", x"00", x"00", 
x"8c", x"84", x"d8", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"98", x"84", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"88", x"84", x"18", x"00", 
x"93", x"65", x"00", x"00", 
x"8c", x"84", x"d8", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"04", 
x"40", x"d0", x"00", x"03", 
x"40", x"f0", x"00", x"02", 
x"41", x"10", x"00", x"01", 
x"07", x"68", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"07", x"64", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"41", x"02", x"00", x"05", 
x"09", x"20", x"00", x"00", 
x"07", x"68", x"48", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"09", x"00", x"00", x"01", 
x"07", x"64", x"40", x"00", 
x"c0", x"7b", x"00", x"00", 
x"41", x"02", x"00", x"05", 
x"09", x"20", x"00", x"01", 
x"07", x"68", x"48", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"09", x"00", x"00", x"02", 
x"07", x"64", x"40", x"00", 
x"c0", x"9b", x"00", x"00", 
x"40", x"82", x"00", x"05", 
x"09", x"00", x"00", x"02", 
x"07", x"64", x"40", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"84", x"28", x"00", 
x"40", x"82", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"20", x"9b", x"00", x"32", 
x"0b", x"60", x"00", x"02", 
x"20", x"9b", x"00", x"03", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"42", x"00", x"04", 
x"47", x"a7", x"ff", x"ff", 
x"c7", x"a4", x"ff", x"fe", 
x"c7", x"a3", x"ff", x"fd", 
x"c7", x"a2", x"ff", x"fc", 
x"47", x"a2", x"ff", x"fb", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"1a", 
x"08", x"40", x"00", x"00", 
x"c0", x"7d", x"ff", x"fc", 
x"c0", x"9d", x"ff", x"fd", 
x"c0", x"bd", x"ff", x"fe", 
x"40", x"7d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"c7", x"a2", x"ff", x"f9", 
x"08", x"43", x"00", x"00", 
x"80", x"43", x"00", x"00", 
x"80", x"64", x"00", x"00", 
x"80", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"91", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"98", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"f9", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"b0", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"a5", x"10", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c5", x"30", x"00", 
x"84", x"c6", x"18", x"00", 
x"9c", x"c6", x"00", x"00", 
x"40", x"c2", x"00", x"04", 
x"08", x"e0", x"00", x"01", 
x"07", x"66", x"38", x"00", 
x"c0", x"fb", x"00", x"00", 
x"ac", x"e6", x"00", x"02", 
x"08", x"c0", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"c0", x"00", x"17", 
x"08", x"c0", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c5", x"30", x"00", 
x"84", x"c6", x"20", x"00", 
x"9c", x"c6", x"00", x"00", 
x"40", x"c2", x"00", x"04", 
x"08", x"e0", x"00", x"02", 
x"07", x"66", x"38", x"00", 
x"c0", x"fb", x"00", x"00", 
x"ac", x"e6", x"00", x"0a", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"e6", x"00", x"00", 
x"a0", x"c7", x"00", x"02", 
x"08", x"c0", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"c0", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"02", 
x"07", x"64", x"30", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"a5", x"18", x"00", 
x"08", x"c0", x"00", x"03", 
x"07", x"64", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c5", x"30", x"00", 
x"84", x"c6", x"10", x"00", 
x"9c", x"c6", x"00", x"00", 
x"40", x"c2", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"fb", x"00", x"00", 
x"ac", x"e6", x"00", x"02", 
x"08", x"c0", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"c0", x"00", x"17", 
x"08", x"c0", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c5", x"30", x"00", 
x"84", x"c6", x"20", x"00", 
x"9c", x"c6", x"00", x"00", 
x"40", x"c2", x"00", x"04", 
x"08", x"e0", x"00", x"02", 
x"07", x"66", x"38", x"00", 
x"c0", x"fb", x"00", x"00", 
x"ac", x"e6", x"00", x"0a", 
x"08", x"c0", x"00", x"03", 
x"07", x"64", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"e6", x"00", x"00", 
x"a0", x"c7", x"00", x"02", 
x"08", x"c0", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"20", x"c0", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"04", 
x"07", x"64", x"30", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"a5", x"20", x"00", 
x"08", x"c0", x"00", x"05", 
x"07", x"64", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"a5", x"20", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"85", x"20", x"00", 
x"84", x"84", x"10", x"00", 
x"9c", x"84", x"00", x"00", 
x"40", x"c2", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"ac", x"44", x"00", x"1a", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"45", x"10", x"00", 
x"84", x"42", x"18", x"00", 
x"9c", x"42", x"00", x"00", 
x"40", x"42", x"00", x"04", 
x"08", x"60", x"00", x"01", 
x"07", x"62", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"0d", 
x"08", x"40", x"00", x"05", 
x"07", x"64", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"a0", x"43", x"00", x"05", 
x"08", x"40", x"00", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"50", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"c4", x"00", x"00", 
x"ac", x"c5", x"00", x"13", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a5", x"10", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"84", x"a5", x"10", x"00", 
x"08", x"a0", x"00", x"03", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"20", x"00", 
x"84", x"a5", x"10", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"08", x"a0", x"00", x"38", 
x"c0", x"c5", x"00", x"00", 
x"a0", x"a6", x"00", x"02", 
x"08", x"a0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"a0", x"00", x"01", 
x"20", x"a0", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c6", x"10", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"e7", x"18", x"00", 
x"84", x"c6", x"38", x"00", 
x"08", x"a0", x"00", x"03", 
x"07", x"63", x"28", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"e7", x"20", x"00", 
x"84", x"c6", x"38", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"c7", x"a5", x"ff", x"fd", 
x"c7", x"a6", x"ff", x"fc", 
x"47", x"a2", x"ff", x"fb", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"05", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"62", x"00", x"01", 
x"0b", x"60", x"00", x"03", 
x"20", x"7b", x"00", x"26", 
x"c0", x"7d", x"ff", x"fc", 
x"8c", x"83", x"18", x"00", 
x"c0", x"bd", x"ff", x"fd", 
x"8c", x"a5", x"10", x"00", 
x"88", x"84", x"28", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"ac", x"82", x"00", x"1c", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"0d", 
x"08", x"40", x"00", x"00", 
x"94", x"84", x"00", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"60", x"00", x"04", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"94", x"84", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"60", x"00", x"04", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"c0", x"7d", x"ff", x"fc", 
x"8c", x"83", x"18", x"00", 
x"c0", x"bd", x"ff", x"fd", 
x"8c", x"a5", x"10", x"00", 
x"88", x"84", x"28", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"ac", x"82", x"00", x"1c", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"0d", 
x"08", x"40", x"00", x"00", 
x"94", x"84", x"00", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"60", x"00", x"04", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"94", x"84", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"60", x"00", x"04", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"04", 
x"40", x"d0", x"00", x"03", 
x"40", x"f0", x"00", x"02", 
x"41", x"10", x"00", x"01", 
x"07", x"68", x"10", x"00", 
x"41", x"1b", x"00", x"00", 
x"09", x"20", x"00", x"00", 
x"07", x"64", x"48", x"00", 
x"c0", x"5b", x"00", x"00", 
x"41", x"28", x"00", x"05", 
x"09", x"40", x"00", x"00", 
x"07", x"69", x"50", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"09", x"20", x"00", x"01", 
x"07", x"64", x"48", x"00", 
x"c0", x"7b", x"00", x"00", 
x"41", x"28", x"00", x"05", 
x"09", x"40", x"00", x"01", 
x"07", x"69", x"50", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"09", x"20", x"00", x"02", 
x"07", x"64", x"48", x"00", 
x"c0", x"9b", x"00", x"00", 
x"40", x"88", x"00", x"05", 
x"09", x"20", x"00", x"02", 
x"07", x"64", x"48", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"84", x"28", x"00", 
x"40", x"83", x"00", x"01", 
x"07", x"64", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"48", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"20", x"5b", x"00", x"0c", 
x"0b", x"60", x"00", x"02", 
x"20", x"5b", x"00", x"05", 
x"08", x"64", x"00", x"00", 
x"08", x"48", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"08", x"48", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"08", x"48", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"50", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"a0", x"00", x"38", 
x"c0", x"65", x"00", x"00", 
x"ac", x"62", x"00", x"0c", 
x"08", x"a0", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"03", 
x"07", x"64", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"07", x"62", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"bb", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"c6", x"00", x"00", 
x"a0", x"a6", x"00", x"02", 
x"08", x"c0", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"c0", x"00", x"01", 
x"20", x"c0", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c6", x"10", x"00", 
x"08", x"c0", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"84", x"c6", x"10", x"00", 
x"08", x"c0", x"00", x"03", 
x"07", x"63", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"42", x"20", x"00", 
x"84", x"c6", x"10", x"00", 
x"08", x"c0", x"00", x"03", 
x"07", x"64", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"66", x"30", x"00", 
x"8c", x"a5", x"10", x"00", 
x"88", x"63", x"28", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"ac", x"62", x"00", x"18", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"0b", 
x"08", x"40", x"00", x"00", 
x"94", x"63", x"00", x"00", 
x"84", x"c6", x"18", x"00", 
x"08", x"80", x"00", x"04", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"c6", x"10", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"94", x"63", x"00", x"00", 
x"88", x"c6", x"18", x"00", 
x"08", x"80", x"00", x"04", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"c6", x"10", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"04", 
x"40", x"b0", x"00", x"03", 
x"40", x"d0", x"00", x"02", 
x"40", x"f0", x"00", x"01", 
x"07", x"67", x"10", x"00", 
x"40", x"fb", x"00", x"00", 
x"41", x"07", x"00", x"0a", 
x"09", x"20", x"00", x"00", 
x"07", x"68", x"48", x"00", 
x"c0", x"5b", x"00", x"00", 
x"09", x"20", x"00", x"01", 
x"07", x"68", x"48", x"00", 
x"c0", x"7b", x"00", x"00", 
x"09", x"20", x"00", x"02", 
x"07", x"68", x"48", x"00", 
x"c0", x"9b", x"00", x"00", 
x"41", x"23", x"00", x"01", 
x"07", x"69", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"41", x"27", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"21", x"3b", x"00", x"0e", 
x"0b", x"60", x"00", x"02", 
x"21", x"3b", x"00", x"06", 
x"08", x"88", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"47", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"08", x"88", x"00", x"00", 
x"08", x"47", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"08", x"82", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"08", x"47", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"80", x"00", x"06", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"60", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"20", x"60", x"00", x"06", 
x"08", x"60", x"00", x"01", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"50", 
x"08", x"60", x"00", x"00", 
x"40", x"bd", x"ff", x"ff", 
x"40", x"c5", x"00", x"06", 
x"08", x"e0", x"00", x"00", 
x"07", x"64", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"e0", x"00", x"38", 
x"c0", x"67", x"00", x"00", 
x"ac", x"62", x"00", x"24", 
x"20", x"c0", x"00", x"12", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"10", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"23", 
x"20", x"c0", x"00", x"11", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"11", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"60", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"20", x"60", x"00", x"06", 
x"08", x"60", x"00", x"03", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"50", 
x"08", x"60", x"00", x"02", 
x"40", x"bd", x"ff", x"ff", 
x"40", x"c5", x"00", x"06", 
x"08", x"e0", x"00", x"01", 
x"07", x"64", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"e0", x"00", x"38", 
x"c0", x"67", x"00", x"00", 
x"ac", x"62", x"00", x"24", 
x"20", x"c0", x"00", x"12", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"01", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"03", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"10", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"01", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"03", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"23", 
x"20", x"c0", x"00", x"11", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"01", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"03", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"20", x"00", x"00", x"11", 
x"40", x"c5", x"00", x"04", 
x"08", x"e0", x"00", x"01", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"03", 
x"08", x"c0", x"00", x"37", 
x"c0", x"46", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"64", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"a0", x"43", x"00", x"02", 
x"08", x"60", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"20", x"60", x"00", x"06", 
x"08", x"60", x"00", x"05", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"04", 
x"40", x"bd", x"ff", x"ff", 
x"40", x"c5", x"00", x"06", 
x"08", x"e0", x"00", x"02", 
x"07", x"64", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"e0", x"00", x"38", 
x"c0", x"67", x"00", x"00", 
x"ac", x"62", x"00", x"24", 
x"20", x"c0", x"00", x"12", 
x"40", x"a5", x"00", x"04", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"05", 
x"08", x"a0", x"00", x"37", 
x"c0", x"45", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"a5", x"00", x"04", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"05", 
x"08", x"a0", x"00", x"37", 
x"c0", x"45", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"20", x"c0", x"00", x"11", 
x"40", x"a5", x"00", x"04", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"05", 
x"08", x"a0", x"00", x"37", 
x"c0", x"45", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"a5", x"00", x"04", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"05", 
x"08", x"a0", x"00", x"37", 
x"c0", x"45", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"04", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"a3", x"00", x"04", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"a3", x"00", x"04", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"83", x"00", x"04", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"64", x"00", x"00", 
x"ac", x"43", x"00", x"02", 
x"08", x"80", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"20", x"80", x"00", x"26", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"36", 
x"c0", x"65", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"40", x"a3", x"00", x"04", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"98", x"63", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"40", x"a3", x"00", x"04", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"98", x"63", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"03", 
x"40", x"63", x"00", x"04", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"98", x"63", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"80", x"00", x"05", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fd", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"05", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"82", x"00", x"04", 
x"08", x"a0", x"00", x"00", 
x"07", x"64", x"28", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"98", x"63", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"40", x"82", x"00", x"04", 
x"08", x"a0", x"00", x"01", 
x"07", x"64", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"84", x"28", x"00", 
x"98", x"84", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"40", x"82", x"00", x"04", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"98", x"a5", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"fd", 
x"07", x"65", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"40", x"82", x"00", x"03", 
x"20", x"80", x"00", x"56", 
x"08", x"80", x"00", x"01", 
x"08", x"c0", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"40", x"c2", x"00", x"09", 
x"08", x"e0", x"00", x"01", 
x"07", x"66", x"38", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"fb", x"00", x"00", 
x"40", x"c2", x"00", x"09", 
x"08", x"e0", x"00", x"02", 
x"07", x"66", x"38", x"00", 
x"c1", x"1b", x"00", x"00", 
x"8c", x"e7", x"40", x"00", 
x"84", x"c6", x"38", x"00", 
x"08", x"c0", x"00", x"31", 
x"c0", x"e6", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"88", x"63", x"30", x"00", 
x"07", x"65", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"08", x"c0", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"c2", x"00", x"09", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"63", x"30", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"db", x"00", x"00", 
x"40", x"c2", x"00", x"09", 
x"08", x"e0", x"00", x"02", 
x"07", x"66", x"38", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"c6", x"38", x"00", 
x"84", x"63", x"30", x"00", 
x"08", x"c0", x"00", x"31", 
x"c0", x"c6", x"00", x"00", 
x"8c", x"63", x"30", x"00", 
x"88", x"84", x"18", x"00", 
x"07", x"65", x"20", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"80", x"00", x"03", 
x"08", x"c0", x"00", x"01", 
x"07", x"63", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"c2", x"00", x"09", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"08", x"c0", x"00", x"00", 
x"07", x"63", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"40", x"42", x"00", x"09", 
x"08", x"60", x"00", x"01", 
x"07", x"62", x"18", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"84", x"30", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"40", x"00", x"31", 
x"c0", x"82", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"88", x"a5", x"18", x"00", 
x"07", x"65", x"20", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"a0", x"43", x"00", x"09", 
x"08", x"40", x"00", x"04", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"65", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"65", x"10", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"07", x"65", x"10", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"a0", x"43", x"00", x"09", 
x"08", x"40", x"00", x"04", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"07", x"65", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"a2", x"00", x"01", 
x"40", x"c2", x"00", x"00", 
x"40", x"e4", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"20", x"fb", x"00", x"2c", 
x"0b", x"60", x"00", x"02", 
x"20", x"fb", x"00", x"15", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a5", x"ff", x"fc", 
x"08", x"64", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0b", x"b6", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a5", x"ff", x"fc", 
x"08", x"64", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0b", x"5c", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a5", x"ff", x"fc", 
x"08", x"64", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"a4", x"00", x"0a", 
x"40", x"c4", x"00", x"01", 
x"08", x"e0", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"07", x"62", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"41", x"04", x"00", x"05", 
x"09", x"20", x"00", x"00", 
x"07", x"68", x"48", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"07", x"65", x"38", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"e0", x"00", x"01", 
x"09", x"00", x"00", x"01", 
x"07", x"62", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"41", x"04", x"00", x"05", 
x"09", x"20", x"00", x"01", 
x"07", x"68", x"48", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"07", x"65", x"38", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"e0", x"00", x"02", 
x"09", x"00", x"00", x"02", 
x"07", x"62", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"41", x"04", x"00", x"05", 
x"09", x"20", x"00", x"02", 
x"07", x"68", x"48", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"07", x"65", x"38", x"00", 
x"c7", x"62", x"00", x"00", 
x"0b", x"60", x"00", x"02", 
x"20", x"db", x"00", x"34", 
x"0b", x"60", x"00", x"02", 
x"2c", x"db", x"00", x"2f", 
x"08", x"e0", x"00", x"00", 
x"07", x"65", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"e0", x"00", x"01", 
x"07", x"65", x"38", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"e0", x"00", x"02", 
x"07", x"65", x"38", x"00", 
x"c0", x"9b", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a5", x"ff", x"fc", 
x"47", x"a6", x"ff", x"fb", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"05", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"03", 
x"40", x"7d", x"ff", x"fb", 
x"0b", x"60", x"00", x"03", 
x"20", x"7b", x"00", x"0a", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"c0", x"00", x"03", 
x"40", x"84", x"00", x"04", 
x"08", x"e0", x"00", x"00", 
x"07", x"65", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"e0", x"00", x"01", 
x"07", x"65", x"38", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"e0", x"00", x"02", 
x"07", x"65", x"38", x"00", 
x"c0", x"9b", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a6", x"ff", x"fa", 
x"47", x"a5", x"ff", x"fc", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"91", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"9c", x"42", x"00", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"ac", x"a2", x"00", x"1a", 
x"9c", x"63", x"00", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"ac", x"43", x"00", x"0e", 
x"9c", x"84", x"00", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"02", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"ac", x"44", x"00", x"02", 
x"40", x"42", x"00", x"06", 
x"33", x"e0", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"07", x"05", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"62", x"00", x"01", 
x"0b", x"60", x"00", x"03", 
x"20", x"7b", x"00", x"0e", 
x"40", x"42", x"00", x"06", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"63", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"40", x"42", x"00", x"06", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"62", x"00", x"05", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"42", x"28", x"00", 
x"40", x"62", x"00", x"05", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"63", x"28", x"00", 
x"40", x"62", x"00", x"05", 
x"08", x"80", x"00", x"02", 
x"07", x"63", x"20", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"84", x"28", x"00", 
x"40", x"62", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"20", x"7b", x"00", x"1a", 
x"0b", x"60", x"00", x"02", 
x"20", x"7b", x"00", x"01", 
x"20", x"00", x"ff", x"c2", 
x"40", x"62", x"00", x"04", 
x"47", x"a2", x"ff", x"ff", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"91", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"42", x"00", x"06", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"ac", x"62", x"00", x"05", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"20", x"00", x"ff", x"84", 
x"40", x"90", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"40", x"bb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"bb", x"00", x"35", 
x"07", x"64", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"c7", x"a4", x"ff", x"fe", 
x"c7", x"a3", x"ff", x"fd", 
x"c7", x"a2", x"ff", x"fc", 
x"47", x"a4", x"ff", x"fb", 
x"47", x"a3", x"ff", x"fa", 
x"47", x"a2", x"ff", x"f9", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0d", x"7e", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f9", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"9b", x"00", x"1a", 
x"40", x"bd", x"ff", x"fb", 
x"07", x"65", x"20", x"00", 
x"40", x"9b", x"00", x"00", 
x"c0", x"5d", x"ff", x"fc", 
x"c0", x"7d", x"ff", x"fd", 
x"c0", x"9d", x"ff", x"fe", 
x"47", x"a2", x"ff", x"f8", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0d", x"7e", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f8", 
x"08", x"42", x"00", x"01", 
x"c0", x"5d", x"ff", x"fc", 
x"c0", x"7d", x"ff", x"fd", 
x"c0", x"9d", x"ff", x"fe", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"ff", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"07", 
x"40", x"b0", x"00", x"06", 
x"40", x"d0", x"00", x"05", 
x"40", x"f0", x"00", x"04", 
x"41", x"10", x"00", x"03", 
x"41", x"30", x"00", x"02", 
x"41", x"50", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"41", x"7b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"21", x"7b", x"00", x"86", 
x"07", x"63", x"10", x"00", 
x"41", x"7b", x"00", x"00", 
x"47", x"aa", x"ff", x"ff", 
x"47", x"a9", x"ff", x"fe", 
x"47", x"a8", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"b0", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"47", x"ab", x"ff", x"f9", 
x"47", x"a6", x"ff", x"f8", 
x"47", x"a5", x"ff", x"f7", 
x"08", x"67", x"00", x"00", 
x"08", x"4b", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"08", x"89", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0e", x"06", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f7", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"20", x"40", x"00", x"07", 
x"08", x"40", x"00", x"30", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"40", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"08", x"40", x"00", x"00", 
x"20", x"40", x"00", x"53", 
x"08", x"40", x"00", x"2f", 
x"c0", x"62", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"10", x"00", 
x"c0", x"9b", x"00", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"84", x"10", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"64", x"10", x"00", 
x"c0", x"bb", x"00", x"00", 
x"84", x"84", x"28", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"63", x"10", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a5", x"10", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"64", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"a5", x"10", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"5b", x"00", x"2e", 
x"40", x"9d", x"ff", x"f8", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"c7", x"a5", x"ff", x"f6", 
x"c7", x"a4", x"ff", x"f5", 
x"c7", x"a3", x"ff", x"f4", 
x"80", x"43", x"00", x"00", 
x"80", x"64", x"00", x"00", 
x"80", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0d", x"7e", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"20", x"40", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"c0", x"5d", x"ff", x"f4", 
x"c0", x"7d", x"ff", x"f5", 
x"c0", x"9d", x"ff", x"f6", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"ff", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0e", x"5b", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f9", 
x"40", x"7d", x"ff", x"f8", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"02", 
x"40", x"b0", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"40", x"db", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"db", x"00", x"1a", 
x"07", x"65", x"30", x"00", 
x"40", x"bb", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fd", 
x"08", x"65", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0e", x"8e", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"05", 
x"40", x"b0", x"00", x"04", 
x"40", x"d0", x"00", x"03", 
x"40", x"f0", x"00", x"02", 
x"41", x"10", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"41", x"3b", x"00", x"00", 
x"09", x"40", x"00", x"00", 
x"07", x"69", x"50", x"00", 
x"41", x"5b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"21", x"5b", x"00", x"69", 
x"0b", x"60", x"00", x"63", 
x"21", x"5b", x"00", x"4f", 
x"47", x"a9", x"ff", x"ff", 
x"47", x"a6", x"ff", x"fe", 
x"47", x"a5", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"b0", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"67", x"00", x"00", 
x"08", x"4a", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"08", x"88", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0e", x"b9", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"36", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"2e", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"28", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0e", x"cc", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"15", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0e", x"d8", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"b0", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"69", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0f", x"05", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"20", x"40", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"09", 
x"40", x"d0", x"00", x"08", 
x"40", x"f0", x"00", x"07", 
x"41", x"10", x"00", x"06", 
x"41", x"30", x"00", x"05", 
x"41", x"50", x"00", x"04", 
x"41", x"70", x"00", x"03", 
x"41", x"90", x"00", x"02", 
x"41", x"b0", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"41", x"db", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"21", x"db", x"00", x"e2", 
x"47", x"ad", x"ff", x"ff", 
x"47", x"aa", x"ff", x"fe", 
x"47", x"ac", x"ff", x"fd", 
x"47", x"ab", x"ff", x"fc", 
x"47", x"a6", x"ff", x"fb", 
x"47", x"a5", x"ff", x"fa", 
x"47", x"a7", x"ff", x"f9", 
x"47", x"a4", x"ff", x"f8", 
x"47", x"a3", x"ff", x"f7", 
x"47", x"b0", x"ff", x"f6", 
x"47", x"a2", x"ff", x"f5", 
x"47", x"ae", x"ff", x"f4", 
x"47", x"a9", x"ff", x"f3", 
x"08", x"64", x"00", x"00", 
x"08", x"4e", x"00", x"00", 
x"0a", x"08", x"00", x"00", 
x"08", x"86", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0f", x"36", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"20", x"40", x"00", x"ba", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"ac", x"43", x"00", x"02", 
x"08", x"60", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"20", x"60", x"00", x"a7", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"60", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"20", x"60", x"00", x"96", 
x"08", x"60", x"00", x"2f", 
x"c0", x"63", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"bd", x"ff", x"f8", 
x"07", x"65", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"dd", x"ff", x"fb", 
x"07", x"66", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"65", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"84", x"10", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"66", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"84", x"84", x"28", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"65", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a5", x"10", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"66", x"18", x"00", 
x"c0", x"db", x"00", x"00", 
x"84", x"a5", x"30", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"dd", x"ff", x"f7", 
x"07", x"66", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"7b", x"00", x"55", 
x"40", x"fd", x"ff", x"f3", 
x"07", x"67", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"47", x"a2", x"ff", x"f2", 
x"c7", x"a2", x"ff", x"f1", 
x"c7", x"a5", x"ff", x"f0", 
x"c7", x"a4", x"ff", x"ef", 
x"c7", x"a3", x"ff", x"ee", 
x"08", x"43", x"00", x"00", 
x"80", x"43", x"00", x"00", 
x"80", x"64", x"00", x"00", 
x"80", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"ed", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0d", x"7e", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"13", 
x"20", x"40", x"00", x"08", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"c0", x"5d", x"ff", x"ee", 
x"c0", x"7d", x"ff", x"ef", 
x"c0", x"9d", x"ff", x"f0", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"ff", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ed", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"0f", x"96", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"13", 
x"20", x"40", x"00", x"24", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"c0", x"5d", x"ff", x"f1", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"c0", x"5d", x"ff", x"ee", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"c0", x"5d", x"ff", x"ef", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"c0", x"5d", x"ff", x"f0", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"f4", 
x"07", x"63", x"10", x"00", 
x"47", x"64", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"f2", 
x"07", x"63", x"10", x"00", 
x"47", x"64", x"00", x"00", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"fd", x"ff", x"f4", 
x"07", x"64", x"18", x"00", 
x"47", x"67", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"08", x"85", x"00", x"00", 
x"0a", x"03", x"00", x"00", 
x"08", x"66", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"40", x"7d", x"ff", x"f3", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"08", 
x"40", x"5d", x"ff", x"f5", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"02", 
x"40", x"d0", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"40", x"fb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"fb", x"00", x"35", 
x"07", x"66", x"38", x"00", 
x"40", x"fb", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a4", x"ff", x"fe", 
x"47", x"a5", x"ff", x"fd", 
x"47", x"a6", x"ff", x"fc", 
x"47", x"a3", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"67", x"00", x"00", 
x"08", x"48", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"1a", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"9b", x"00", x"1a", 
x"40", x"bd", x"ff", x"fc", 
x"07", x"65", x"20", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"40", x"dd", x"ff", x"fe", 
x"40", x"fd", x"ff", x"fd", 
x"47", x"a2", x"ff", x"f9", 
x"08", x"64", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"08", x"86", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"33", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"5d", x"ff", x"f9", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fe", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"07", 
x"40", x"d0", x"00", x"06", 
x"40", x"f0", x"00", x"05", 
x"41", x"10", x"00", x"04", 
x"41", x"30", x"00", x"03", 
x"41", x"50", x"00", x"02", 
x"41", x"70", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"41", x"9b", x"00", x"00", 
x"09", x"a0", x"00", x"00", 
x"07", x"6c", x"68", x"00", 
x"41", x"bb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"21", x"bb", x"00", x"93", 
x"0b", x"60", x"00", x"63", 
x"21", x"bb", x"00", x"62", 
x"47", x"a9", x"ff", x"ff", 
x"47", x"aa", x"ff", x"fe", 
x"47", x"ab", x"ff", x"fd", 
x"47", x"ac", x"ff", x"fc", 
x"47", x"a5", x"ff", x"fb", 
x"47", x"a7", x"ff", x"fa", 
x"47", x"a4", x"ff", x"f9", 
x"47", x"a3", x"ff", x"f8", 
x"47", x"b0", x"ff", x"f7", 
x"47", x"a2", x"ff", x"f6", 
x"08", x"64", x"00", x"00", 
x"08", x"4d", x"00", x"00", 
x"0a", x"08", x"00", x"00", 
x"08", x"86", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"62", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"20", x"40", x"00", x"44", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"33", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"5b", x"00", x"25", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"f9", 
x"40", x"dd", x"ff", x"fe", 
x"08", x"62", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"08", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"83", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"8f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"6c", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"bb", x"00", x"27", 
x"07", x"6b", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"47", x"a3", x"ff", x"f8", 
x"47", x"b0", x"ff", x"f7", 
x"47", x"a2", x"ff", x"f6", 
x"47", x"a4", x"ff", x"f9", 
x"47", x"ac", x"ff", x"fc", 
x"47", x"a9", x"ff", x"ff", 
x"08", x"65", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0a", x"0a", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"c7", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"d3", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"42", x"00", x"01", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"03", 
x"40", x"90", x"00", x"02", 
x"40", x"b0", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"08", x"e0", x"00", x"2d", 
x"c0", x"47", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"08", x"e0", x"00", x"00", 
x"07", x"65", x"38", x"00", 
x"40", x"bb", x"00", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"08", x"82", x"00", x"00", 
x"0a", x"03", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"10", x"f7", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"2e", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"07", 
x"08", x"40", x"00", x"2c", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"09", 
x"40", x"d0", x"00", x"08", 
x"40", x"f0", x"00", x"07", 
x"41", x"10", x"00", x"06", 
x"41", x"30", x"00", x"05", 
x"41", x"50", x"00", x"04", 
x"41", x"70", x"00", x"03", 
x"41", x"90", x"00", x"02", 
x"41", x"b0", x"00", x"01", 
x"41", x"c4", x"00", x"00", 
x"07", x"63", x"10", x"00", 
x"41", x"fb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"21", x"fb", x"00", x"e2", 
x"47", x"ad", x"ff", x"ff", 
x"47", x"aa", x"ff", x"fe", 
x"47", x"ac", x"ff", x"fd", 
x"47", x"ab", x"ff", x"fc", 
x"47", x"a6", x"ff", x"fb", 
x"47", x"ae", x"ff", x"fa", 
x"47", x"a5", x"ff", x"f9", 
x"47", x"a8", x"ff", x"f8", 
x"47", x"a4", x"ff", x"f7", 
x"47", x"a3", x"ff", x"f6", 
x"47", x"b0", x"ff", x"f5", 
x"47", x"a2", x"ff", x"f4", 
x"47", x"af", x"ff", x"f3", 
x"47", x"a9", x"ff", x"f2", 
x"08", x"64", x"00", x"00", 
x"08", x"4f", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"11", x"2d", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"20", x"40", x"00", x"ba", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f8", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"63", x"00", x"00", 
x"ac", x"43", x"00", x"02", 
x"08", x"60", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"20", x"60", x"00", x"a7", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"60", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"20", x"60", x"00", x"96", 
x"08", x"60", x"00", x"2f", 
x"c0", x"63", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"07", x"65", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"dd", x"ff", x"fb", 
x"07", x"66", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"65", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"84", x"10", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"66", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"84", x"84", x"28", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"65", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a5", x"10", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"66", x"18", x"00", 
x"c0", x"db", x"00", x"00", 
x"84", x"a5", x"30", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"bd", x"ff", x"f6", 
x"07", x"65", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"7b", x"00", x"55", 
x"40", x"dd", x"ff", x"f2", 
x"07", x"66", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"47", x"a2", x"ff", x"f1", 
x"c7", x"a2", x"ff", x"f0", 
x"c7", x"a5", x"ff", x"ef", 
x"c7", x"a4", x"ff", x"ee", 
x"c7", x"a3", x"ff", x"ed", 
x"08", x"43", x"00", x"00", 
x"80", x"43", x"00", x"00", 
x"80", x"64", x"00", x"00", 
x"80", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"0d", x"7e", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"20", x"40", x"00", x"08", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"bd", x"ff", x"f5", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"c0", x"5d", x"ff", x"ed", 
x"c0", x"7d", x"ff", x"ee", 
x"c0", x"9d", x"ff", x"ef", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"ff", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"11", x"8d", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"20", x"40", x"00", x"24", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"f9", 
x"c0", x"5d", x"ff", x"f0", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"c0", x"5d", x"ff", x"ed", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"c0", x"5d", x"ff", x"ee", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"c0", x"5d", x"ff", x"ef", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"63", x"10", x"00", 
x"47", x"64", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"f1", 
x"07", x"63", x"10", x"00", 
x"47", x"64", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"bd", x"ff", x"f5", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"bd", x"ff", x"f5", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"dd", x"ff", x"f3", 
x"07", x"64", x"18", x"00", 
x"47", x"66", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f5", 
x"0a", x"03", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"bd", x"ff", x"f5", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"bd", x"ff", x"f5", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"f2", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"20", x"40", x"00", x"08", 
x"40", x"5d", x"ff", x"f4", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f7", 
x"40", x"bd", x"ff", x"f5", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"02", 
x"40", x"d0", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"40", x"fb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"fb", x"00", x"35", 
x"07", x"66", x"38", x"00", 
x"40", x"fb", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a4", x"ff", x"fe", 
x"47", x"a5", x"ff", x"fd", 
x"47", x"a6", x"ff", x"fc", 
x"47", x"a3", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"67", x"00", x"00", 
x"08", x"48", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"11", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"9b", x"00", x"1a", 
x"40", x"bd", x"ff", x"fc", 
x"07", x"65", x"20", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"40", x"dd", x"ff", x"fe", 
x"40", x"fd", x"ff", x"fd", 
x"47", x"a2", x"ff", x"f9", 
x"08", x"64", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"08", x"86", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"2a", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"5d", x"ff", x"f9", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fe", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"06", 
x"40", x"d0", x"00", x"05", 
x"40", x"f0", x"00", x"04", 
x"41", x"10", x"00", x"03", 
x"41", x"30", x"00", x"02", 
x"41", x"50", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"41", x"7b", x"00", x"00", 
x"09", x"80", x"00", x"00", 
x"07", x"6b", x"60", x"00", 
x"41", x"9b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"21", x"9b", x"00", x"92", 
x"0b", x"60", x"00", x"63", 
x"21", x"9b", x"00", x"61", 
x"47", x"a8", x"ff", x"ff", 
x"47", x"a9", x"ff", x"fe", 
x"47", x"aa", x"ff", x"fd", 
x"47", x"ab", x"ff", x"fc", 
x"47", x"a5", x"ff", x"fb", 
x"47", x"a7", x"ff", x"fa", 
x"47", x"a4", x"ff", x"f9", 
x"47", x"a3", x"ff", x"f8", 
x"47", x"b0", x"ff", x"f7", 
x"47", x"a2", x"ff", x"f6", 
x"08", x"64", x"00", x"00", 
x"08", x"4c", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"57", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"20", x"40", x"00", x"44", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"ac", x"62", x"00", x"33", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"5b", x"00", x"25", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"f9", 
x"40", x"dd", x"ff", x"fe", 
x"08", x"62", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"08", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"78", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"84", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"6b", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"0b", x"60", x"ff", x"ff", 
x"20", x"bb", x"00", x"27", 
x"07", x"6a", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"47", x"a3", x"ff", x"f8", 
x"47", x"b0", x"ff", x"f7", 
x"47", x"a2", x"ff", x"f6", 
x"47", x"a4", x"ff", x"f9", 
x"47", x"ab", x"ff", x"fc", 
x"47", x"a8", x"ff", x"ff", 
x"08", x"65", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0a", x"09", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"bc", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"c8", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f6", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f7", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"42", x"00", x"01", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"03", 
x"40", x"90", x"00", x"02", 
x"40", x"b0", x"00", x"01", 
x"08", x"c0", x"00", x"00", 
x"08", x"e0", x"00", x"2d", 
x"c0", x"47", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"08", x"e0", x"00", x"00", 
x"07", x"65", x"38", x"00", 
x"40", x"bb", x"00", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"08", x"82", x"00", x"00", 
x"0a", x"03", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"12", x"ec", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"2e", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"07", 
x"08", x"40", x"00", x"2c", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"02", 
x"40", x"90", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"07", x"64", x"28", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a4", x"ff", x"ff", 
x"08", x"84", x"ff", x"ff", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"a0", x"43", x"00", x"0d", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"05", 
x"08", x"40", x"00", x"36", 
x"c0", x"42", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"37", 
x"c0", x"42", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"40", x"a2", x"00", x"04", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"40", x"a2", x"00", x"04", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"40", x"42", x"00", x"04", 
x"08", x"a0", x"00", x"02", 
x"07", x"62", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"02", 
x"40", x"90", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"07", x"64", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"a2", x"00", x"05", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"64", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"a2", x"00", x"05", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"9b", x"00", x"00", 
x"40", x"82", x"00", x"05", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"84", x"28", x"00", 
x"40", x"82", x"00", x"04", 
x"08", x"a0", x"00", x"00", 
x"07", x"64", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a2", x"28", x"00", 
x"40", x"82", x"00", x"04", 
x"08", x"a0", x"00", x"01", 
x"07", x"64", x"28", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c3", x"30", x"00", 
x"40", x"82", x"00", x"04", 
x"08", x"a0", x"00", x"02", 
x"07", x"64", x"28", x"00", 
x"c0", x"fb", x"00", x"00", 
x"8c", x"e4", x"38", x"00", 
x"40", x"82", x"00", x"03", 
x"20", x"80", x"00", x"3b", 
x"08", x"80", x"00", x"00", 
x"40", x"a2", x"00", x"09", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c1", x"1b", x"00", x"00", 
x"8d", x"03", x"40", x"00", 
x"40", x"a2", x"00", x"09", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c1", x"3b", x"00", x"00", 
x"8d", x"24", x"48", x"00", 
x"85", x"08", x"48", x"00", 
x"08", x"a0", x"00", x"31", 
x"c1", x"25", x"00", x"00", 
x"8d", x"08", x"48", x"00", 
x"84", x"a5", x"40", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"40", x"a2", x"00", x"09", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"a2", x"28", x"00", 
x"40", x"a2", x"00", x"09", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c1", x"1b", x"00", x"00", 
x"8c", x"84", x"40", x"00", 
x"84", x"a5", x"20", x"00", 
x"08", x"a0", x"00", x"31", 
x"c0", x"85", x"00", x"00", 
x"8c", x"a5", x"20", x"00", 
x"84", x"c6", x"28", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"40", x"a2", x"00", x"09", 
x"08", x"c0", x"00", x"01", 
x"07", x"65", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"42", x"20", x"00", 
x"40", x"a2", x"00", x"09", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"84", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"31", 
x"c0", x"65", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"84", x"e7", x"10", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"67", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"20", x"00", x"ec", x"6f", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"07", x"63", x"20", x"00", 
x"c7", x"67", x"00", x"00", 
x"40", x"42", x"00", x"06", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"20", x"00", x"ec", x"61", 
x"40", x"90", x"00", x"01", 
x"40", x"a2", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"40", x"e2", x"00", x"08", 
x"09", x"00", x"00", x"00", 
x"07", x"67", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"c0", x"00", x"01", 
x"40", x"e2", x"00", x"08", 
x"09", x"00", x"00", x"01", 
x"07", x"67", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"c0", x"00", x"02", 
x"40", x"e2", x"00", x"08", 
x"09", x"00", x"00", x"02", 
x"07", x"67", x"40", x"00", 
x"c0", x"5b", x"00", x"00", 
x"07", x"64", x"30", x"00", 
x"c7", x"62", x"00", x"00", 
x"0b", x"60", x"00", x"01", 
x"20", x"bb", x"01", x"0e", 
x"0b", x"60", x"00", x"02", 
x"20", x"bb", x"00", x"ee", 
x"0b", x"60", x"00", x"03", 
x"20", x"bb", x"00", x"b7", 
x"0b", x"60", x"00", x"04", 
x"20", x"bb", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"a2", x"00", x"05", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"40", x"a2", x"00", x"04", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"94", x"63", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"a2", x"00", x"05", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"40", x"a2", x"00", x"04", 
x"08", x"c0", x"00", x"02", 
x"07", x"65", x"30", x"00", 
x"c0", x"9b", x"00", x"00", 
x"94", x"84", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"8c", x"82", x"10", x"00", 
x"8c", x"a3", x"18", x"00", 
x"84", x"84", x"28", x"00", 
x"9c", x"a2", x"00", x"00", 
x"08", x"a0", x"00", x"2b", 
x"c0", x"c5", x"00", x"00", 
x"ac", x"c5", x"00", x"02", 
x"08", x"a0", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"c7", x"a4", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"20", x"a0", x"00", x"03", 
x"08", x"a0", x"00", x"2a", 
x"c0", x"45", x"00", x"00", 
x"20", x"00", x"00", x"0f", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"9c", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"13", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"08", x"40", x"00", x"29", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"40", x"00", x"28", 
x"c0", x"62", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"b8", x"62", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"40", x"62", x"00", x"05", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"40", x"42", x"00", x"04", 
x"08", x"60", x"00", x"01", 
x"07", x"62", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"94", x"84", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"c0", x"9d", x"ff", x"fe", 
x"9c", x"a4", x"00", x"00", 
x"08", x"40", x"00", x"2b", 
x"c0", x"c2", x"00", x"00", 
x"ac", x"c5", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"40", x"00", x"00", 
x"20", x"40", x"00", x"26", 
x"08", x"40", x"00", x"2a", 
x"c0", x"62", x"00", x"00", 
x"b8", x"83", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"40", x"00", x"27", 
x"c0", x"82", x"00", x"00", 
x"08", x"40", x"00", x"31", 
x"c0", x"a2", x"00", x"00", 
x"88", x"a5", x"10", x"00", 
x"8c", x"a5", x"28", x"00", 
x"88", x"84", x"28", x"00", 
x"08", x"40", x"00", x"31", 
x"c0", x"42", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"8c", x"42", x"10", x"00", 
x"88", x"84", x"10", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"ac", x"44", x"00", x"07", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"26", 
x"c0", x"43", x"00", x"00", 
x"8c", x"42", x"20", x"00", 
x"08", x"60", x"00", x"25", 
x"c0", x"63", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"93", x"64", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"9c", x"63", x"00", x"00", 
x"c7", x"a2", x"ff", x"fb", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"13", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"40", x"00", x"29", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"40", x"00", x"28", 
x"c0", x"62", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"b8", x"62", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"27", 
x"c0", x"62", x"00", x"00", 
x"08", x"40", x"00", x"31", 
x"c0", x"82", x"00", x"00", 
x"c0", x"bd", x"ff", x"fb", 
x"88", x"84", x"28", x"00", 
x"8c", x"84", x"20", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"40", x"00", x"31", 
x"c0", x"82", x"00", x"00", 
x"88", x"84", x"10", x"00", 
x"8c", x"84", x"20", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"ac", x"43", x"00", x"07", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"26", 
x"c0", x"43", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"60", x"00", x"25", 
x"c0", x"63", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"a2", x"00", x"05", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"7b", x"00", x"00", 
x"40", x"42", x"00", x"05", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"8c", x"42", x"10", x"00", 
x"8c", x"63", x"18", x"00", 
x"84", x"42", x"18", x"00", 
x"94", x"42", x"00", x"00", 
x"08", x"40", x"00", x"24", 
x"c0", x"62", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"b8", x"62", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"28", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"8c", x"42", x"10", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"26", 
x"c0", x"63", x"00", x"00", 
x"8c", x"62", x"18", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"80", x"00", x"37", 
x"c0", x"64", x"00", x"00", 
x"88", x"63", x"10", x"00", 
x"08", x"80", x"00", x"26", 
x"c0", x"44", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"40", x"00", x"23", 
x"c0", x"62", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"8c", x"42", x"10", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"26", 
x"c0", x"63", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"80", x"00", x"26", 
x"c0", x"64", x"00", x"00", 
x"08", x"80", x"00", x"37", 
x"c0", x"84", x"00", x"00", 
x"88", x"84", x"10", x"00", 
x"8c", x"63", x"20", x"00", 
x"07", x"63", x"10", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"a2", x"00", x"05", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"22", 
x"c0", x"65", x"00", x"00", 
x"8c", x"62", x"18", x"00", 
x"b8", x"63", x"00", x"00", 
x"08", x"a0", x"00", x"21", 
x"c0", x"85", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"a0", x"00", x"24", 
x"c0", x"65", x"00", x"00", 
x"ac", x"62", x"00", x"1f", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"05", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"22", 
x"c0", x"62", x"00", x"00", 
x"8c", x"62", x"18", x"00", 
x"b8", x"63", x"00", x"00", 
x"08", x"40", x"00", x"21", 
x"c0", x"82", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"24", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"06", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"26", 
x"c0", x"43", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c0", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"05", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"22", 
x"c0", x"62", x"00", x"00", 
x"8c", x"62", x"18", x"00", 
x"b8", x"63", x"00", x"00", 
x"08", x"40", x"00", x"21", 
x"c0", x"82", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"40", x"00", x"24", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"06", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"26", 
x"c0", x"43", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"02", 
x"40", x"50", x"00", x"01", 
x"08", x"80", x"00", x"38", 
x"c0", x"a4", x"00", x"00", 
x"ac", x"45", x"00", x"02", 
x"08", x"80", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"20", x"80", x"00", x"28", 
x"47", x"a2", x"ff", x"ff", 
x"c7", x"a4", x"ff", x"fe", 
x"c7", x"a3", x"ff", x"fd", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"a0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"fd", 
x"ac", x"62", x"00", x"1b", 
x"8c", x"63", x"18", x"00", 
x"8c", x"63", x"18", x"00", 
x"c0", x"5d", x"ff", x"fe", 
x"8c", x"63", x"10", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"ff", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"ac", x"62", x"00", x"19", 
x"8c", x"63", x"18", x"00", 
x"8c", x"63", x"18", x"00", 
x"8c", x"63", x"20", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"02", 
x"07", x"62", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"08", 
x"40", x"b0", x"00", x"07", 
x"40", x"d0", x"00", x"06", 
x"40", x"f0", x"00", x"05", 
x"41", x"10", x"00", x"04", 
x"41", x"30", x"00", x"03", 
x"41", x"50", x"00", x"02", 
x"41", x"70", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"65", x"10", x"00", 
x"40", x"bb", x"00", x"00", 
x"41", x"85", x"00", x"01", 
x"47", x"ab", x"ff", x"ff", 
x"47", x"a7", x"ff", x"fe", 
x"47", x"ac", x"ff", x"fd", 
x"47", x"a4", x"ff", x"fc", 
x"47", x"a6", x"ff", x"fb", 
x"47", x"a5", x"ff", x"fa", 
x"47", x"a9", x"ff", x"f9", 
x"47", x"aa", x"ff", x"f8", 
x"c7", x"a3", x"ff", x"f7", 
x"c7", x"a2", x"ff", x"f6", 
x"47", x"a3", x"ff", x"f5", 
x"47", x"b0", x"ff", x"f4", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"4c", x"00", x"00", 
x"0a", x"08", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"15", x"9d", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"20", x"40", x"00", x"5d", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"f8", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"14", x"42", x"00", x"02", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"83", x"00", x"00", 
x"20", x"44", x"00", x"09", 
x"40", x"5d", x"ff", x"f3", 
x"08", x"42", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"f6", 
x"c0", x"7d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f5", 
x"40", x"9d", x"ff", x"f4", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"fb", 
x"07", x"65", x"20", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"bd", x"ff", x"fc", 
x"08", x"64", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"15", x"c3", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"20", x"40", x"00", x"09", 
x"40", x"5d", x"ff", x"f3", 
x"08", x"42", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"f6", 
x"c0", x"7d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f5", 
x"40", x"9d", x"ff", x"f4", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"40", x"62", x"00", x"00", 
x"40", x"9d", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"fa", 
x"c0", x"62", x"00", x"02", 
x"c0", x"9d", x"ff", x"f6", 
x"8c", x"a3", x"20", x"00", 
x"8c", x"a5", x"10", x"00", 
x"40", x"5d", x"ff", x"fd", 
x"40", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f5", 
x"c7", x"a5", x"ff", x"f2", 
x"c7", x"a3", x"ff", x"f1", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"c0", x"7d", x"ff", x"f1", 
x"8c", x"63", x"10", x"00", 
x"c0", x"5d", x"ff", x"f2", 
x"c0", x"9d", x"ff", x"f7", 
x"40", x"5d", x"ff", x"ff", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"15", x"f2", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"40", x"5d", x"ff", x"f3", 
x"08", x"42", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"f6", 
x"c0", x"7d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f5", 
x"40", x"9d", x"ff", x"f4", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f3", 
x"08", x"42", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"f6", 
x"c0", x"7d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f5", 
x"40", x"9d", x"ff", x"f4", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"b0", x"00", x"18", 
x"40", x"d0", x"00", x"17", 
x"40", x"f0", x"00", x"16", 
x"41", x"10", x"00", x"15", 
x"41", x"30", x"00", x"14", 
x"41", x"50", x"00", x"13", 
x"41", x"70", x"00", x"12", 
x"41", x"90", x"00", x"11", 
x"41", x"b0", x"00", x"10", 
x"41", x"d0", x"00", x"0f", 
x"41", x"f0", x"00", x"0e", 
x"47", x"a7", x"ff", x"ff", 
x"40", x"f0", x"00", x"0d", 
x"47", x"a6", x"ff", x"fe", 
x"40", x"d0", x"00", x"0c", 
x"47", x"a6", x"ff", x"fd", 
x"40", x"d0", x"00", x"0b", 
x"47", x"ac", x"ff", x"fc", 
x"41", x"90", x"00", x"0a", 
x"47", x"a6", x"ff", x"fb", 
x"40", x"d0", x"00", x"09", 
x"47", x"a9", x"ff", x"fa", 
x"41", x"30", x"00", x"08", 
x"47", x"ab", x"ff", x"f9", 
x"41", x"70", x"00", x"07", 
x"47", x"ae", x"ff", x"f8", 
x"41", x"d0", x"00", x"06", 
x"47", x"a7", x"ff", x"f7", 
x"40", x"f0", x"00", x"05", 
x"47", x"a8", x"ff", x"f6", 
x"41", x"10", x"00", x"04", 
x"47", x"a9", x"ff", x"f5", 
x"41", x"30", x"00", x"03", 
x"47", x"a5", x"ff", x"f4", 
x"40", x"b0", x"00", x"02", 
x"47", x"ab", x"ff", x"f3", 
x"41", x"70", x"00", x"01", 
x"0b", x"60", x"00", x"04", 
x"2c", x"5b", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"47", x"ab", x"ff", x"f2", 
x"41", x"64", x"00", x"02", 
x"47", x"b0", x"ff", x"f1", 
x"c7", x"a3", x"ff", x"f0", 
x"47", x"a4", x"ff", x"ef", 
x"47", x"aa", x"ff", x"ee", 
x"47", x"a7", x"ff", x"ed", 
x"47", x"a9", x"ff", x"ec", 
x"47", x"a8", x"ff", x"eb", 
x"47", x"af", x"ff", x"ea", 
x"47", x"ae", x"ff", x"e9", 
x"47", x"ad", x"ff", x"e8", 
x"47", x"a5", x"ff", x"e7", 
x"c7", x"a2", x"ff", x"e6", 
x"47", x"ac", x"ff", x"e5", 
x"47", x"a3", x"ff", x"e4", 
x"47", x"a2", x"ff", x"e3", 
x"47", x"ab", x"ff", x"e2", 
x"08", x"43", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"e1", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"16", x"47", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1f", 
x"20", x"40", x"01", x"52", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"e9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"ea", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"83", x"00", x"02", 
x"40", x"a3", x"00", x"07", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"c0", x"7d", x"ff", x"e6", 
x"8c", x"42", x"18", x"00", 
x"40", x"a3", x"00", x"01", 
x"47", x"a4", x"ff", x"e1", 
x"c7", x"a2", x"ff", x"e0", 
x"47", x"a2", x"ff", x"df", 
x"47", x"a3", x"ff", x"de", 
x"0b", x"60", x"00", x"01", 
x"20", x"bb", x"00", x"18", 
x"0b", x"60", x"00", x"02", 
x"20", x"bb", x"00", x"0b", 
x"40", x"bd", x"ff", x"ed", 
x"08", x"43", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"16", x"69", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"20", x"00", x"00", x"0a", 
x"40", x"bd", x"ff", x"ec", 
x"08", x"43", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"16", x"74", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"20", x"00", x"00", x"0b", 
x"40", x"bd", x"ff", x"e4", 
x"40", x"dd", x"ff", x"eb", 
x"08", x"45", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"16", x"80", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"40", x"5d", x"ff", x"ee", 
x"40", x"7d", x"ff", x"f3", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"40", x"5d", x"ff", x"de", 
x"40", x"7d", x"ff", x"f3", 
x"40", x"9d", x"ff", x"f4", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"16", x"92", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"40", x"5d", x"ff", x"df", 
x"14", x"42", x"00", x"02", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f5", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"40", x"7d", x"ff", x"e3", 
x"40", x"9d", x"ff", x"e2", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"ef", 
x"40", x"a2", x"00", x"01", 
x"07", x"65", x"18", x"00", 
x"40", x"bb", x"00", x"00", 
x"40", x"dd", x"ff", x"f3", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"40", x"5d", x"ff", x"ef", 
x"40", x"62", x"00", x"03", 
x"40", x"9d", x"ff", x"de", 
x"40", x"a4", x"00", x"07", 
x"08", x"c0", x"00", x"00", 
x"07", x"65", x"30", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"a0", x"00", x"31", 
x"c0", x"65", x"00", x"00", 
x"ac", x"62", x"00", x"02", 
x"08", x"a0", x"00", x"01", 
x"20", x"00", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"20", x"a0", x"00", x"05", 
x"08", x"a0", x"00", x"00", 
x"40", x"dd", x"ff", x"e3", 
x"07", x"63", x"30", x"00", 
x"47", x"65", x"00", x"00", 
x"20", x"00", x"00", x"2b", 
x"08", x"a0", x"00", x"01", 
x"40", x"dd", x"ff", x"e3", 
x"07", x"63", x"30", x"00", 
x"47", x"65", x"00", x"00", 
x"40", x"62", x"00", x"04", 
x"07", x"63", x"30", x"00", 
x"40", x"bb", x"00", x"00", 
x"40", x"fd", x"ff", x"f6", 
x"47", x"a3", x"ff", x"dd", 
x"08", x"67", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"dc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"24", 
x"40", x"5d", x"ff", x"e3", 
x"40", x"7d", x"ff", x"dd", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"80", x"00", x"20", 
x"c0", x"44", x"00", x"00", 
x"c0", x"7d", x"ff", x"e0", 
x"8c", x"42", x"18", x"00", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"dc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"e1", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"24", 
x"40", x"5d", x"ff", x"ef", 
x"40", x"62", x"00", x"07", 
x"40", x"9d", x"ff", x"e3", 
x"07", x"63", x"20", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"f7", 
x"08", x"43", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"0b", x"bd", x"ff", x"dc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"24", 
x"08", x"40", x"00", x"1f", 
x"c0", x"42", x"00", x"00", 
x"40", x"5d", x"ff", x"e4", 
x"40", x"7d", x"ff", x"f7", 
x"c7", x"a2", x"ff", x"dc", 
x"0b", x"bd", x"ff", x"db", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"25", 
x"c0", x"7d", x"ff", x"dc", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"e4", 
x"40", x"7d", x"ff", x"f7", 
x"0b", x"bd", x"ff", x"db", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"a0", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"25", 
x"40", x"5d", x"ff", x"de", 
x"40", x"62", x"00", x"07", 
x"08", x"80", x"00", x"01", 
x"07", x"63", x"20", x"00", 
x"c0", x"5b", x"00", x"00", 
x"c0", x"7d", x"ff", x"e6", 
x"8c", x"43", x"10", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"f8", 
x"07", x"65", x"20", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"bd", x"ff", x"f9", 
x"c7", x"a2", x"ff", x"db", 
x"08", x"43", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"da", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"17", x"12", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"26", 
x"20", x"40", x"00", x"01", 
x"20", x"00", x"00", x"1e", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"e5", 
x"0b", x"bd", x"ff", x"da", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"26", 
x"98", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"e0", 
x"8c", x"42", x"18", x"00", 
x"40", x"5d", x"ff", x"e4", 
x"40", x"7d", x"ff", x"e5", 
x"c7", x"a2", x"ff", x"da", 
x"0b", x"bd", x"ff", x"d9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"27", 
x"98", x"62", x"00", x"00", 
x"c0", x"5d", x"ff", x"da", 
x"c0", x"9d", x"ff", x"db", 
x"40", x"5d", x"ff", x"f2", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"d9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"17", x"32", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"27", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"f3", 
x"0b", x"bd", x"ff", x"d9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"27", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"9d", x"ff", x"fc", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"d9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"17", x"48", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"27", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fd", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"e0", 
x"c0", x"7d", x"ff", x"db", 
x"40", x"7d", x"ff", x"e4", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"d9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"17", x"59", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"27", 
x"08", x"40", x"00", x"1e", 
x"c0", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"e6", 
x"ac", x"62", x"00", x"3c", 
x"40", x"5d", x"ff", x"e3", 
x"0b", x"60", x"00", x"04", 
x"2f", x"62", x"00", x"1f", 
x"08", x"62", x"00", x"01", 
x"08", x"80", x"ff", x"ff", 
x"40", x"bd", x"ff", x"e2", 
x"07", x"65", x"18", x"00", 
x"47", x"64", x"00", x"00", 
x"40", x"7d", x"ff", x"e1", 
x"0b", x"60", x"00", x"02", 
x"20", x"7b", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"de", 
x"40", x"63", x"00", x"07", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"42", x"20", x"00", 
x"8c", x"43", x"10", x"00", 
x"08", x"42", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"ff", 
x"07", x"64", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c0", x"9d", x"ff", x"f0", 
x"84", x"64", x"18", x"00", 
x"40", x"7d", x"ff", x"e4", 
x"40", x"9d", x"ff", x"ef", 
x"40", x"bd", x"ff", x"f1", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"7d", x"ff", x"e1", 
x"0b", x"60", x"00", x"02", 
x"20", x"7b", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"de", 
x"40", x"63", x"00", x"07", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"42", x"20", x"00", 
x"8c", x"43", x"10", x"00", 
x"08", x"42", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"ff", 
x"07", x"64", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"c0", x"9d", x"ff", x"f0", 
x"84", x"64", x"18", x"00", 
x"40", x"7d", x"ff", x"e4", 
x"40", x"9d", x"ff", x"ef", 
x"40", x"bd", x"ff", x"f1", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"ff", x"ff", 
x"40", x"7d", x"ff", x"e3", 
x"40", x"9d", x"ff", x"e2", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"20", x"60", x"00", x"2c", 
x"40", x"5d", x"ff", x"e4", 
x"40", x"7d", x"ff", x"e5", 
x"0b", x"bd", x"ff", x"d9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"27", 
x"98", x"42", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"20", 
x"8c", x"62", x"10", x"00", 
x"8c", x"63", x"10", x"00", 
x"c0", x"5d", x"ff", x"e6", 
x"8c", x"63", x"10", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"e7", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"63", x"10", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"e8", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"02", 
x"07", x"64", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"07", x"64", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"0e", 
x"40", x"90", x"00", x"0d", 
x"40", x"b0", x"00", x"0c", 
x"40", x"d0", x"00", x"0b", 
x"40", x"f0", x"00", x"0a", 
x"41", x"10", x"00", x"09", 
x"41", x"30", x"00", x"08", 
x"41", x"50", x"00", x"07", 
x"41", x"70", x"00", x"06", 
x"41", x"90", x"00", x"05", 
x"41", x"b0", x"00", x"04", 
x"41", x"d0", x"00", x"03", 
x"41", x"f0", x"00", x"02", 
x"47", x"ad", x"ff", x"ff", 
x"41", x"b0", x"00", x"01", 
x"47", x"af", x"ff", x"fe", 
x"47", x"a4", x"ff", x"fd", 
x"47", x"ad", x"ff", x"fc", 
x"c7", x"a2", x"ff", x"fb", 
x"47", x"a9", x"ff", x"fa", 
x"47", x"a8", x"ff", x"f9", 
x"47", x"a5", x"ff", x"f8", 
x"47", x"a6", x"ff", x"f7", 
x"47", x"ab", x"ff", x"f6", 
x"47", x"a3", x"ff", x"f5", 
x"47", x"ae", x"ff", x"f4", 
x"47", x"a2", x"ff", x"f3", 
x"47", x"a7", x"ff", x"f2", 
x"47", x"ac", x"ff", x"f1", 
x"0a", x"0a", x"00", x"00", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"17", x"f2", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"20", x"40", x"00", x"e7", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"f1", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"f2", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"f3", 
x"40", x"63", x"00", x"00", 
x"40", x"82", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"20", x"9b", x"00", x"92", 
x"0b", x"60", x"00", x"02", 
x"20", x"9b", x"00", x"48", 
x"40", x"7d", x"ff", x"ff", 
x"47", x"a2", x"ff", x"f0", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"0b", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f5", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"16", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f7", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f8", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"24", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"20", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f9", 
x"40", x"7d", x"ff", x"fa", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"98", x"42", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"0b", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"42", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"7d", x"ff", x"fd", 
x"20", x"00", x"e8", x"62", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"42", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"7d", x"ff", x"fd", 
x"20", x"00", x"e8", x"55", 
x"40", x"7d", x"ff", x"fe", 
x"47", x"a2", x"ff", x"f0", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"53", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f5", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"5e", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f7", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f8", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"6c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"20", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f9", 
x"40", x"7d", x"ff", x"fa", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"98", x"42", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"0b", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"42", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"7d", x"ff", x"fd", 
x"20", x"00", x"e8", x"1a", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"42", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"7d", x"ff", x"fd", 
x"20", x"00", x"e8", x"0d", 
x"40", x"9d", x"ff", x"f4", 
x"47", x"a2", x"ff", x"f0", 
x"08", x"43", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"9c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"7d", x"ff", x"f6", 
x"40", x"9d", x"ff", x"f5", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"a7", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f7", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f8", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"18", x"b5", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"20", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f9", 
x"40", x"7d", x"ff", x"fa", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"98", x"42", x"00", x"00", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"43", x"00", x"0b", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"42", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"7d", x"ff", x"fd", 
x"20", x"00", x"e7", x"d1", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"c0", x"7d", x"ff", x"fb", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"f0", 
x"40", x"42", x"00", x"07", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"8c", x"43", x"10", x"00", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"7d", x"ff", x"fd", 
x"20", x"00", x"e7", x"c4", 
x"33", x"e0", x"00", x"00", 
x"40", x"d0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"65", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"62", x"28", x"00", 
x"40", x"fb", x"00", x"00", 
x"40", x"e7", x"00", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"47", x"b0", x"ff", x"fd", 
x"47", x"a6", x"ff", x"fc", 
x"47", x"a5", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"47", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"40", x"00", x"38", 
x"c0", x"62", x"00", x"00", 
x"ac", x"62", x"00", x"1c", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"62", x"00", x"01", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"a0", x"00", x"1d", 
x"c0", x"65", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"40", x"bd", x"ff", x"fc", 
x"08", x"43", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"04", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"a2", x"ff", x"fe", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"ff", 
x"40", x"dd", x"ff", x"fd", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"1c", 
x"c0", x"65", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"40", x"bd", x"ff", x"fc", 
x"08", x"44", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"1f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"a2", x"ff", x"fe", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"ff", 
x"40", x"dd", x"ff", x"fd", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"b0", x"00", x"05", 
x"40", x"d0", x"00", x"04", 
x"40", x"f0", x"00", x"03", 
x"41", x"10", x"00", x"02", 
x"41", x"30", x"00", x"01", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a8", x"ff", x"fe", 
x"47", x"a6", x"ff", x"fd", 
x"47", x"a7", x"ff", x"fc", 
x"47", x"a4", x"ff", x"fb", 
x"47", x"a5", x"ff", x"fa", 
x"47", x"a9", x"ff", x"f9", 
x"47", x"a2", x"ff", x"f8", 
x"20", x"40", x"00", x"2a", 
x"09", x"40", x"00", x"00", 
x"07", x"69", x"50", x"00", 
x"41", x"5b", x"00", x"00", 
x"47", x"aa", x"ff", x"f7", 
x"08", x"64", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"52", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"5f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"20", x"00", x"00", x"00", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"01", 
x"20", x"5b", x"01", x"5a", 
x"08", x"60", x"00", x"01", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f6", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"82", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f6", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"8f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"02", 
x"20", x"5b", x"00", x"ac", 
x"08", x"60", x"00", x"02", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f5", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0c", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f4", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"b1", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0c", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f5", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f4", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"be", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0c", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"03", 
x"20", x"5b", x"00", x"55", 
x"08", x"60", x"00", x"03", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f4", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"e0", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f4", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"19", x"ed", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"0d", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"35", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"03", 
x"20", x"5b", x"00", x"55", 
x"08", x"60", x"00", x"03", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f4", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"5f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f4", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"6c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"8c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"b4", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"02", 
x"20", x"5b", x"00", x"ac", 
x"08", x"60", x"00", x"02", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f5", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"de", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f5", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1a", x"eb", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"03", 
x"20", x"5b", x"00", x"55", 
x"08", x"60", x"00", x"03", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f4", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"0d", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f4", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"1a", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"3a", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"62", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"03", 
x"20", x"5b", x"00", x"55", 
x"08", x"60", x"00", x"03", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"fb", 
x"47", x"a3", x"ff", x"f4", 
x"08", x"66", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fd", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"8c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f4", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"99", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f8", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"b9", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"04", 
x"20", x"5b", x"00", x"25", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f9", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1b", x"e1", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"f3", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"dd", x"ff", x"fe", 
x"0a", x"06", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"03", 
x"40", x"b0", x"00", x"02", 
x"40", x"d0", x"00", x"01", 
x"40", x"e2", x"00", x"05", 
x"41", x"02", x"00", x"07", 
x"41", x"22", x"00", x"01", 
x"41", x"42", x"00", x"04", 
x"07", x"67", x"18", x"00", 
x"40", x"fb", x"00", x"00", 
x"47", x"a6", x"ff", x"ff", 
x"47", x"a5", x"ff", x"fe", 
x"47", x"aa", x"ff", x"fd", 
x"47", x"a4", x"ff", x"fc", 
x"47", x"a9", x"ff", x"fb", 
x"47", x"a3", x"ff", x"fa", 
x"47", x"a8", x"ff", x"f9", 
x"47", x"a2", x"ff", x"f8", 
x"08", x"67", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"42", x"00", x"06", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"18", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"bd", x"ff", x"fb", 
x"07", x"65", x"18", x"00", 
x"40", x"bb", x"00", x"00", 
x"40", x"dd", x"ff", x"fc", 
x"08", x"64", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"08", x"85", x"00", x"00", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1c", x"19", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"fd", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"5d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"ff", 
x"20", x"00", x"e4", x"d5", 
x"40", x"f0", x"00", x"02", 
x"41", x"10", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"05", 
x"09", x"22", x"ff", x"ff", 
x"07", x"64", x"48", x"00", 
x"41", x"3b", x"00", x"00", 
x"41", x"29", x"00", x"05", 
x"07", x"64", x"10", x"00", 
x"41", x"5b", x"00", x"00", 
x"41", x"4a", x"00", x"05", 
x"09", x"62", x"00", x"01", 
x"07", x"64", x"58", x"00", 
x"41", x"7b", x"00", x"00", 
x"41", x"6b", x"00", x"05", 
x"07", x"65", x"10", x"00", 
x"40", x"bb", x"00", x"00", 
x"40", x"a5", x"00", x"05", 
x"07", x"63", x"30", x"00", 
x"40", x"7b", x"00", x"00", 
x"47", x"a7", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"47", x"a4", x"ff", x"fd", 
x"47", x"a5", x"ff", x"fc", 
x"47", x"ab", x"ff", x"fb", 
x"47", x"aa", x"ff", x"fa", 
x"47", x"a8", x"ff", x"f9", 
x"47", x"a6", x"ff", x"f8", 
x"47", x"a9", x"ff", x"f7", 
x"08", x"48", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"f7", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"c2", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"c2", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"fb", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"c2", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"c2", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"40", x"5d", x"ff", x"fe", 
x"40", x"7d", x"ff", x"fd", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"04", 
x"40", x"7d", x"ff", x"f8", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"f9", 
x"20", x"00", x"e4", x"7a", 
x"40", x"90", x"00", x"01", 
x"0b", x"60", x"00", x"04", 
x"2c", x"7b", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"a2", x"00", x"02", 
x"07", x"65", x"18", x"00", 
x"40", x"bb", x"00", x"00", 
x"0b", x"60", x"00", x"00", 
x"2f", x"65", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"a2", x"00", x"03", 
x"07", x"65", x"18", x"00", 
x"40", x"bb", x"00", x"00", 
x"20", x"a0", x"00", x"12", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"b0", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1c", x"94", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"63", x"00", x"01", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"08", x"a0", x"00", x"01", 
x"07", x"64", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"08", x"c3", x"00", x"01", 
x"2c", x"a6", x"00", x"11", 
x"0b", x"60", x"00", x"00", 
x"2c", x"7b", x"00", x"0d", 
x"08", x"60", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"82", x"00", x"01", 
x"2c", x"64", x"00", x"06", 
x"0b", x"60", x"00", x"00", 
x"2c", x"5b", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"07", x"64", x"10", x"00", 
x"40", x"fb", x"00", x"00", 
x"40", x"e7", x"00", x"02", 
x"07", x"67", x"30", x"00", 
x"40", x"fb", x"00", x"00", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"40", x"7b", x"00", x"00", 
x"20", x"67", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"07", x"65", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"40", x"7b", x"00", x"00", 
x"20", x"67", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"02", 
x"07", x"63", x"30", x"00", 
x"40", x"7b", x"00", x"00", 
x"20", x"67", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"42", x"00", x"01", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"02", 
x"07", x"62", x"30", x"00", 
x"40", x"5b", x"00", x"00", 
x"20", x"47", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"41", x"10", x"00", x"02", 
x"41", x"30", x"00", x"01", 
x"07", x"65", x"10", x"00", 
x"41", x"5b", x"00", x"00", 
x"0b", x"60", x"00", x"04", 
x"2c", x"fb", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"41", x"6a", x"00", x"02", 
x"07", x"6b", x"38", x"00", 
x"41", x"7b", x"00", x"00", 
x"0b", x"60", x"00", x"00", 
x"2f", x"6b", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"47", x"a9", x"ff", x"ff", 
x"47", x"a6", x"ff", x"fe", 
x"47", x"a4", x"ff", x"fd", 
x"47", x"a3", x"ff", x"fc", 
x"47", x"b0", x"ff", x"fb", 
x"47", x"aa", x"ff", x"fa", 
x"47", x"a7", x"ff", x"f9", 
x"47", x"a8", x"ff", x"f8", 
x"47", x"a2", x"ff", x"f7", 
x"47", x"a5", x"ff", x"f6", 
x"08", x"64", x"00", x"00", 
x"08", x"85", x"00", x"00", 
x"08", x"a6", x"00", x"00", 
x"08", x"c7", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"1c", x"b9", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"20", x"40", x"00", x"28", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"42", x"00", x"03", 
x"40", x"dd", x"ff", x"f9", 
x"07", x"62", x"30", x"00", 
x"40", x"5b", x"00", x"00", 
x"20", x"40", x"00", x"18", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"f6", 
x"40", x"bd", x"ff", x"fe", 
x"40", x"fd", x"ff", x"ff", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1d", x"14", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f9", 
x"08", x"e2", x"00", x"01", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"bd", x"ff", x"f6", 
x"40", x"dd", x"ff", x"fe", 
x"41", x"1d", x"ff", x"fb", 
x"0a", x"08", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"e6", x"00", x"01", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"bd", x"ff", x"f6", 
x"40", x"dd", x"ff", x"fe", 
x"41", x"1d", x"ff", x"fb", 
x"0a", x"08", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f6", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"7d", x"ff", x"f9", 
x"40", x"9d", x"ff", x"f8", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"50", x"00", x"01", 
x"08", x"60", x"00", x"50", 
x"47", x"a2", x"ff", x"ff", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"33", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"20", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"20", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"f6", 
x"40", x"50", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c0", x"5b", x"00", x"00", 
x"b0", x"62", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"0b", x"60", x"00", x"ff", 
x"2c", x"7b", x"00", x"08", 
x"08", x"60", x"00", x"ff", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"20", x"00", x"00", x"10", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"08", 
x"08", x"60", x"00", x"00", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"20", x"00", x"00", x"06", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"20", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"01", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"b0", x"42", x"00", x"00", 
x"0b", x"60", x"00", x"ff", 
x"2c", x"5b", x"00", x"2c", 
x"08", x"40", x"00", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"20", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"b0", x"42", x"00", x"00", 
x"0b", x"60", x"00", x"ff", 
x"2c", x"5b", x"00", x"08", 
x"08", x"40", x"00", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"ae", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"08", 
x"08", x"40", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"a4", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"9d", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"2c", 
x"08", x"40", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"20", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"b0", x"42", x"00", x"00", 
x"0b", x"60", x"00", x"ff", 
x"2c", x"5b", x"00", x"08", 
x"08", x"40", x"00", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"80", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"08", 
x"08", x"40", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"76", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"6f", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"20", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"65", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"02", 
x"40", x"7d", x"ff", x"ff", 
x"07", x"63", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"b0", x"42", x"00", x"00", 
x"0b", x"60", x"00", x"ff", 
x"2c", x"5b", x"00", x"08", 
x"08", x"40", x"00", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"55", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"08", 
x"08", x"40", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"4b", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"67", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"40", x"00", x"0a", 
x"20", x"00", x"0c", x"44", 
x"40", x"90", x"00", x"06", 
x"40", x"b0", x"00", x"05", 
x"40", x"d0", x"00", x"04", 
x"40", x"f0", x"00", x"03", 
x"41", x"10", x"00", x"02", 
x"41", x"30", x"00", x"01", 
x"0b", x"60", x"00", x"04", 
x"2c", x"7b", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"41", x"42", x"00", x"02", 
x"07", x"6a", x"18", x"00", 
x"41", x"5b", x"00", x"00", 
x"0b", x"60", x"00", x"00", 
x"2f", x"6a", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"41", x"42", x"00", x"03", 
x"07", x"6a", x"18", x"00", 
x"41", x"5b", x"00", x"00", 
x"21", x"40", x"00", x"58", 
x"41", x"42", x"00", x"06", 
x"09", x"60", x"00", x"00", 
x"07", x"6a", x"58", x"00", 
x"41", x"5b", x"00", x"00", 
x"09", x"60", x"00", x"38", 
x"c0", x"4b", x"00", x"00", 
x"09", x"60", x"00", x"00", 
x"07", x"69", x"58", x"00", 
x"c7", x"62", x"00", x"00", 
x"09", x"60", x"00", x"01", 
x"07", x"69", x"58", x"00", 
x"c7", x"62", x"00", x"00", 
x"09", x"60", x"00", x"02", 
x"07", x"69", x"58", x"00", 
x"c7", x"62", x"00", x"00", 
x"41", x"62", x"00", x"07", 
x"41", x"82", x"00", x"01", 
x"07", x"68", x"50", x"00", 
x"41", x"1b", x"00", x"00", 
x"07", x"6b", x"18", x"00", 
x"41", x"5b", x"00", x"00", 
x"07", x"6c", x"18", x"00", 
x"41", x"7b", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a9", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a2", x"ff", x"fc", 
x"47", x"aa", x"ff", x"fb", 
x"47", x"a8", x"ff", x"fa", 
x"47", x"a7", x"ff", x"f9", 
x"47", x"ab", x"ff", x"f8", 
x"47", x"a5", x"ff", x"f7", 
x"47", x"a6", x"ff", x"f6", 
x"08", x"6b", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"f6", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f7", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1e", x"69", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"a0", x"00", x"76", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"7d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"f8", 
x"40", x"dd", x"ff", x"f9", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1e", x"76", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"62", x"00", x"05", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"63", x"20", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"bd", x"ff", x"fe", 
x"08", x"43", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"ff", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"63", x"00", x"01", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"b0", x"00", x"09", 
x"40", x"d0", x"00", x"08", 
x"40", x"f0", x"00", x"07", 
x"41", x"10", x"00", x"06", 
x"41", x"30", x"00", x"05", 
x"41", x"50", x"00", x"04", 
x"41", x"70", x"00", x"03", 
x"41", x"90", x"00", x"02", 
x"41", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"09", x"c0", x"00", x"00", 
x"07", x"69", x"70", x"00", 
x"c0", x"bb", x"00", x"00", 
x"09", x"20", x"00", x"00", 
x"07", x"6d", x"48", x"00", 
x"41", x"3b", x"00", x"00", 
x"11", x"23", x"48", x"00", 
x"b4", x"c9", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"09", x"20", x"00", x"00", 
x"09", x"a0", x"00", x"00", 
x"07", x"68", x"68", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c5", x"30", x"00", 
x"84", x"c6", x"10", x"00", 
x"07", x"6b", x"48", x"00", 
x"c7", x"66", x"00", x"00", 
x"09", x"20", x"00", x"01", 
x"09", x"a0", x"00", x"01", 
x"07", x"68", x"68", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"c5", x"30", x"00", 
x"84", x"c6", x"18", x"00", 
x"07", x"6b", x"48", x"00", 
x"c7", x"66", x"00", x"00", 
x"09", x"20", x"00", x"02", 
x"09", x"a0", x"00", x"02", 
x"07", x"68", x"68", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"84", x"a5", x"20", x"00", 
x"07", x"6b", x"48", x"00", 
x"c7", x"65", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"c7", x"a4", x"ff", x"ff", 
x"c7", x"a3", x"ff", x"fe", 
x"c7", x"a2", x"ff", x"fd", 
x"47", x"b0", x"ff", x"fc", 
x"47", x"ac", x"ff", x"fb", 
x"47", x"a4", x"ff", x"fa", 
x"47", x"ab", x"ff", x"f9", 
x"47", x"a6", x"ff", x"f8", 
x"47", x"a3", x"ff", x"f7", 
x"47", x"a2", x"ff", x"f6", 
x"47", x"a5", x"ff", x"f5", 
x"47", x"a7", x"ff", x"f4", 
x"47", x"aa", x"ff", x"f3", 
x"08", x"68", x"00", x"00", 
x"08", x"4b", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"16", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"38", 
x"c0", x"42", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"f3", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"01", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"63", x"10", x"00", 
x"c7", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f4", 
x"40", x"9d", x"ff", x"f5", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"40", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"f7", 
x"40", x"9d", x"ff", x"f6", 
x"07", x"64", x"18", x"00", 
x"40", x"bb", x"00", x"00", 
x"08", x"c0", x"00", x"38", 
x"c0", x"66", x"00", x"00", 
x"40", x"dd", x"ff", x"f9", 
x"40", x"fd", x"ff", x"f8", 
x"08", x"85", x"00", x"00", 
x"08", x"66", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1e", x"f8", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f6", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"84", x"00", x"00", 
x"40", x"bd", x"ff", x"f3", 
x"08", x"65", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f6", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"40", x"84", x"00", x"06", 
x"08", x"a0", x"00", x"00", 
x"40", x"dd", x"ff", x"fa", 
x"07", x"64", x"28", x"00", 
x"47", x"66", x"00", x"00", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"40", x"fd", x"ff", x"fb", 
x"08", x"65", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"1c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"40", x"5d", x"ff", x"f7", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"82", x"00", x"01", 
x"0b", x"60", x"00", x"05", 
x"2f", x"64", x"00", x"08", 
x"c0", x"5d", x"ff", x"fd", 
x"c0", x"7d", x"ff", x"fe", 
x"c0", x"9d", x"ff", x"ff", 
x"40", x"5d", x"ff", x"f6", 
x"40", x"bd", x"ff", x"fc", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"84", x"ff", x"fb", 
x"c0", x"5d", x"ff", x"fd", 
x"c0", x"7d", x"ff", x"fe", 
x"c0", x"9d", x"ff", x"ff", 
x"40", x"5d", x"ff", x"f6", 
x"40", x"bd", x"ff", x"fc", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"b0", x"00", x"06", 
x"40", x"d0", x"00", x"05", 
x"40", x"f0", x"00", x"04", 
x"41", x"10", x"00", x"03", 
x"41", x"30", x"00", x"02", 
x"41", x"50", x"00", x"01", 
x"09", x"60", x"00", x"00", 
x"07", x"67", x"58", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"e0", x"00", x"01", 
x"07", x"6a", x"38", x"00", 
x"40", x"fb", x"00", x"00", 
x"10", x"63", x"38", x"00", 
x"b4", x"63", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"66", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"8c", x"62", x"18", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"65", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"84", x"63", x"20", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"66", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"82", x"20", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"65", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"84", x"84", x"28", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"66", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"42", x"28", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"65", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"84", x"42", x"28", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"69", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"0a", x"08", x"00", x"00", 
x"83", x"64", x"00", x"00", 
x"80", x"82", x"00", x"00", 
x"80", x"43", x"00", x"00", 
x"80", x"7b", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"f0", x"00", x"06", 
x"41", x"10", x"00", x"05", 
x"41", x"30", x"00", x"04", 
x"41", x"50", x"00", x"03", 
x"41", x"70", x"00", x"02", 
x"41", x"90", x"00", x"01", 
x"09", x"a0", x"00", x"00", 
x"07", x"6b", x"68", x"00", 
x"41", x"7b", x"00", x"00", 
x"2d", x"62", x"00", x"66", 
x"07", x"65", x"10", x"00", 
x"41", x"7b", x"00", x"00", 
x"41", x"6b", x"00", x"00", 
x"47", x"a8", x"ff", x"ff", 
x"47", x"a4", x"ff", x"fe", 
x"47", x"b0", x"ff", x"fd", 
x"47", x"a7", x"ff", x"fc", 
x"47", x"ac", x"ff", x"fb", 
x"47", x"a5", x"ff", x"fa", 
x"47", x"a6", x"ff", x"f9", 
x"47", x"a3", x"ff", x"f8", 
x"47", x"a2", x"ff", x"f7", 
x"47", x"aa", x"ff", x"f6", 
x"08", x"6b", x"00", x"00", 
x"08", x"49", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f9", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"8f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"20", x"40", x"00", x"22", 
x"08", x"e0", x"00", x"00", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"fe", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"f9", 
x"41", x"1d", x"ff", x"ff", 
x"0a", x"08", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"9f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"fc", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"a8", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f7", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"fe", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"f9", 
x"40", x"fd", x"ff", x"fd", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"40", x"dd", x"ff", x"fb", 
x"08", x"65", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"c2", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"fc", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"cb", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"f7", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"fe", 
x"40", x"bd", x"ff", x"fa", 
x"40", x"dd", x"ff", x"f9", 
x"40", x"fd", x"ff", x"fd", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"f0", x"00", x"03", 
x"41", x"10", x"00", x"02", 
x"41", x"30", x"00", x"01", 
x"09", x"40", x"00", x"01", 
x"07", x"69", x"50", x"00", 
x"41", x"5b", x"00", x"00", 
x"2d", x"42", x"00", x"64", 
x"09", x"40", x"00", x"01", 
x"07", x"69", x"50", x"00", 
x"41", x"3b", x"00", x"00", 
x"09", x"29", x"ff", x"ff", 
x"2d", x"22", x"00", x"36", 
x"09", x"22", x"00", x"01", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a6", x"ff", x"fe", 
x"47", x"a5", x"ff", x"fd", 
x"47", x"a4", x"ff", x"fc", 
x"47", x"a3", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"47", x"a7", x"ff", x"f9", 
x"08", x"86", x"00", x"00", 
x"08", x"69", x"00", x"00", 
x"08", x"45", x"00", x"00", 
x"0a", x"08", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"1f", x"f5", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"fc", 
x"40", x"dd", x"ff", x"fd", 
x"40", x"fd", x"ff", x"f9", 
x"0a", x"07", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"20", x"03", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fe", 
x"08", x"c3", x"00", x"02", 
x"0b", x"60", x"00", x"05", 
x"2f", x"66", x"00", x"07", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"bd", x"ff", x"fb", 
x"40", x"fd", x"ff", x"ff", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"c6", x"ff", x"fb", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"bd", x"ff", x"fb", 
x"40", x"fd", x"ff", x"ff", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"47", x"a3", x"ff", x"fb", 
x"47", x"a5", x"ff", x"fd", 
x"47", x"a4", x"ff", x"fc", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a6", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"c5", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"08", x"a4", x"00", x"00", 
x"08", x"83", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"48", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"20", x"2c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"00", x"01", 
x"40", x"7d", x"ff", x"fe", 
x"08", x"c3", x"00", x"02", 
x"0b", x"60", x"00", x"05", 
x"2f", x"66", x"00", x"07", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"bd", x"ff", x"fb", 
x"40", x"fd", x"ff", x"ff", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"c6", x"ff", x"fb", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fd", 
x"40", x"bd", x"ff", x"fb", 
x"40", x"fd", x"ff", x"ff", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"05", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"03", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"40", x"00", x"02", 
x"08", x"60", x"00", x"03", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a2", x"ff", x"fd", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"60", x"00", x"03", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a2", x"ff", x"fc", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"40", x"7d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"40", x"00", x"04", 
x"08", x"60", x"00", x"03", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a2", x"ff", x"fb", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"40", x"7d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"47", x"a2", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"44", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"60", x"00", x"05", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"60", x"00", x"05", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"fd", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"47", x"a2", x"ff", x"fc", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"44", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"47", x"a2", x"ff", x"fb", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"44", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"47", x"a2", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"44", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"08", 
x"44", x"62", x"00", x"07", 
x"40", x"5d", x"ff", x"f9", 
x"44", x"62", x"00", x"06", 
x"40", x"5d", x"ff", x"fa", 
x"44", x"62", x"00", x"05", 
x"40", x"5d", x"ff", x"fb", 
x"44", x"62", x"00", x"04", 
x"40", x"5d", x"ff", x"fc", 
x"44", x"62", x"00", x"03", 
x"40", x"5d", x"ff", x"fd", 
x"44", x"62", x"00", x"02", 
x"40", x"5d", x"ff", x"fe", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"ff", 
x"44", x"62", x"00", x"00", 
x"08", x"43", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"47", x"a3", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"92", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"40", x"7d", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"02", 
x"08", x"44", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"47", x"a3", x"ff", x"fd", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"92", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fe", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"08", x"44", x"00", x"00", 
x"20", x"00", x"ff", x"e0", 
x"40", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"05", 
x"2f", x"62", x"00", x"5d", 
x"8c", x"63", x"18", x"00", 
x"08", x"a0", x"00", x"1e", 
x"c0", x"45", x"00", x"00", 
x"84", x"63", x"10", x"00", 
x"94", x"63", x"00", x"00", 
x"08", x"a0", x"00", x"37", 
x"c0", x"45", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"47", x"a4", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"47", x"b0", x"ff", x"fd", 
x"c7", x"a5", x"ff", x"fc", 
x"47", x"a2", x"ff", x"fb", 
x"c7", x"a3", x"ff", x"fa", 
x"c7", x"a4", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"13", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"c0", x"7d", x"ff", x"f9", 
x"8c", x"42", x"18", x"00", 
x"c7", x"a2", x"ff", x"f8", 
x"0b", x"bd", x"ff", x"f7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"09", 
x"c0", x"7d", x"ff", x"f8", 
x"c7", x"a2", x"ff", x"f7", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"c0", x"7d", x"ff", x"f7", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"c0", x"5d", x"ff", x"fa", 
x"8c", x"63", x"10", x"00", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"42", x"00", x"01", 
x"8c", x"43", x"18", x"00", 
x"08", x"60", x"00", x"1e", 
x"c0", x"83", x"00", x"00", 
x"84", x"42", x"20", x"00", 
x"94", x"42", x"00", x"00", 
x"08", x"60", x"00", x"37", 
x"c0", x"83", x"00", x"00", 
x"93", x"62", x"00", x"00", 
x"8c", x"84", x"d8", x"00", 
x"c7", x"a3", x"ff", x"f6", 
x"47", x"a2", x"ff", x"f5", 
x"c7", x"a2", x"ff", x"f4", 
x"80", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"13", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"c0", x"7d", x"ff", x"fc", 
x"8c", x"42", x"18", x"00", 
x"c7", x"a2", x"ff", x"f3", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"ce", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"c0", x"7d", x"ff", x"f3", 
x"c7", x"a2", x"ff", x"f2", 
x"80", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"9a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"c0", x"7d", x"ff", x"f2", 
x"93", x"62", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"c0", x"5d", x"ff", x"f4", 
x"8c", x"63", x"10", x"00", 
x"c0", x"5d", x"ff", x"f6", 
x"c0", x"9d", x"ff", x"f9", 
x"c0", x"bd", x"ff", x"fc", 
x"40", x"5d", x"ff", x"f5", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"ff", 
x"40", x"bd", x"ff", x"fd", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"8c", x"82", x"10", x"00", 
x"8c", x"a3", x"18", x"00", 
x"84", x"84", x"28", x"00", 
x"08", x"40", x"00", x"37", 
x"c0", x"a2", x"00", x"00", 
x"84", x"84", x"28", x"00", 
x"94", x"84", x"00", x"00", 
x"93", x"64", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"93", x"64", x"00", x"00", 
x"8c", x"63", x"d8", x"00", 
x"08", x"40", x"00", x"37", 
x"c0", x"a2", x"00", x"00", 
x"93", x"64", x"00", x"00", 
x"8c", x"a5", x"d8", x"00", 
x"07", x"65", x"18", x"00", 
x"40", x"5b", x"00", x"00", 
x"07", x"62", x"20", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"64", x"00", x"28", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"98", x"83", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"64", x"00", x"50", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"98", x"82", x"00", x"00", 
x"98", x"c3", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"64", x"00", x"01", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"98", x"82", x"00", x"00", 
x"98", x"c3", x"00", x"00", 
x"98", x"e5", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c7", x"67", x"00", x"00", 
x"08", x"64", x"00", x"29", 
x"07", x"62", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"40", x"63", x"00", x"00", 
x"98", x"82", x"00", x"00", 
x"98", x"c5", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"07", x"63", x"28", x"00", 
x"c7", x"64", x"00", x"00", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c7", x"66", x"00", x"00", 
x"08", x"a0", x"00", x"02", 
x"07", x"63", x"28", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"84", x"00", x"51", 
x"07", x"62", x"20", x"00", 
x"40", x"5b", x"00", x"00", 
x"40", x"42", x"00", x"00", 
x"98", x"a5", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"c7", x"65", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"62", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c7", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"b4", x"62", x"00", x"00", 
x"08", x"c0", x"00", x"1b", 
x"c0", x"86", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"08", x"c0", x"00", x"1a", 
x"c0", x"86", x"00", x"00", 
x"88", x"83", x"20", x"00", 
x"08", x"c0", x"00", x"00", 
x"08", x"e0", x"00", x"38", 
x"c0", x"67", x"00", x"00", 
x"08", x"e0", x"00", x"38", 
x"c0", x"a7", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"c7", x"a2", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a5", x"ff", x"fc", 
x"47", x"a4", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"46", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"83", x"65", x"00", x"00", 
x"80", x"a2", x"00", x"00", 
x"80", x"43", x"00", x"00", 
x"80", x"7b", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"21", x"ec", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"b4", x"42", x"00", x"00", 
x"08", x"60", x"00", x"1b", 
x"c0", x"63", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"60", x"00", x"1e", 
x"c0", x"63", x"00", x"00", 
x"84", x"82", x"18", x"00", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"64", x"00", x"00", 
x"40", x"9d", x"ff", x"fb", 
x"08", x"a4", x"00", x"02", 
x"c0", x"bd", x"ff", x"fe", 
x"40", x"dd", x"ff", x"fd", 
x"40", x"fd", x"ff", x"fc", 
x"08", x"85", x"00", x"00", 
x"08", x"43", x"00", x"00", 
x"0a", x"07", x"00", x"00", 
x"08", x"66", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"22", x"09", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"ff", x"ff", 
x"40", x"7d", x"ff", x"fd", 
x"08", x"63", x"00", x"01", 
x"0b", x"60", x"00", x"05", 
x"2f", x"63", x"00", x"06", 
x"c0", x"5d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"63", x"ff", x"fb", 
x"c0", x"5d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"fb", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"b4", x"42", x"00", x"00", 
x"08", x"c0", x"00", x"1b", 
x"c0", x"66", x"00", x"00", 
x"8c", x"42", x"18", x"00", 
x"08", x"c0", x"00", x"1a", 
x"c0", x"66", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"c0", x"00", x"04", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a4", x"ff", x"fe", 
x"47", x"a3", x"ff", x"fd", 
x"47", x"a2", x"ff", x"fc", 
x"08", x"46", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"22", x"35", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"40", x"5d", x"ff", x"fc", 
x"08", x"42", x"ff", x"ff", 
x"40", x"7d", x"ff", x"fd", 
x"08", x"63", x"00", x"02", 
x"0b", x"60", x"00", x"05", 
x"2f", x"63", x"00", x"06", 
x"40", x"9d", x"ff", x"fe", 
x"08", x"84", x"00", x"04", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"63", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fe", 
x"08", x"84", x"00", x"04", 
x"40", x"bd", x"ff", x"ff", 
x"0a", x"05", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"90", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"a0", x"00", x"03", 
x"08", x"c0", x"00", x"38", 
x"c0", x"46", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fd", 
x"47", x"a4", x"ff", x"fc", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"fb", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"fb", 
x"44", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"10", x"00", 
x"47", x"63", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"60", x"00", x"03", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"f9", 
x"44", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fa", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"10", x"00", 
x"47", x"63", x"00", x"00", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"0a", x"02", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"70", x"00", x"03", 
x"40", x"90", x"00", x"02", 
x"40", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"08", x"c0", x"00", x"78", 
x"08", x"e0", x"00", x"03", 
x"09", x"00", x"00", x"38", 
x"c0", x"48", x"00", x"00", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a5", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fd", 
x"47", x"a4", x"ff", x"fc", 
x"47", x"a6", x"ff", x"fb", 
x"47", x"a3", x"ff", x"fa", 
x"08", x"47", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"f9", 
x"44", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fb", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"40", x"7d", x"ff", x"fd", 
x"40", x"9d", x"ff", x"fc", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"07", x"64", x"18", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"80", x"00", x"76", 
x"08", x"a0", x"00", x"03", 
x"08", x"c0", x"00", x"38", 
x"c0", x"46", x"00", x"00", 
x"47", x"a4", x"ff", x"f8", 
x"47", x"a2", x"ff", x"f7", 
x"08", x"45", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"f6", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"f6", 
x"44", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"9d", x"ff", x"f7", 
x"07", x"64", x"10", x"00", 
x"47", x"63", x"00", x"00", 
x"08", x"60", x"00", x"75", 
x"40", x"5d", x"ff", x"fe", 
x"0a", x"02", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"22", x"f2", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"42", x"ff", x"ff", 
x"40", x"7d", x"ff", x"ff", 
x"0a", x"03", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"90", x"00", x"02", 
x"40", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"63", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"62", x"18", x"00", 
x"40", x"db", x"00", x"00", 
x"08", x"e0", x"00", x"00", 
x"07", x"64", x"38", x"00", 
x"40", x"fb", x"00", x"00", 
x"08", x"e7", x"ff", x"ff", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a5", x"ff", x"fe", 
x"47", x"a4", x"ff", x"fd", 
x"47", x"a2", x"ff", x"fc", 
x"47", x"a3", x"ff", x"fb", 
x"08", x"67", x"00", x"00", 
x"08", x"46", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"23", x"12", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"42", x"ff", x"ff", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"7d", x"ff", x"fc", 
x"07", x"63", x"10", x"00", 
x"40", x"9b", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"40", x"dd", x"ff", x"fd", 
x"07", x"66", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"08", x"a5", x"ff", x"ff", 
x"40", x"dd", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"65", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0a", x"06", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"23", x"2b", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"62", x"ff", x"ff", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"ff", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"70", x"00", x"04", 
x"40", x"90", x"00", x"03", 
x"40", x"b0", x"00", x"02", 
x"40", x"d0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"66", x"10", x"00", 
x"40", x"fb", x"00", x"00", 
x"09", x"00", x"00", x"77", 
x"07", x"67", x"40", x"00", 
x"41", x"1b", x"00", x"00", 
x"09", x"20", x"00", x"00", 
x"07", x"63", x"48", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"63", x"ff", x"ff", 
x"47", x"b0", x"ff", x"ff", 
x"47", x"a6", x"ff", x"fe", 
x"47", x"a2", x"ff", x"fd", 
x"47", x"a7", x"ff", x"fc", 
x"47", x"a5", x"ff", x"fb", 
x"08", x"48", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"23", x"50", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"60", x"00", x"76", 
x"40", x"5d", x"ff", x"fc", 
x"40", x"9d", x"ff", x"fb", 
x"0a", x"04", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"23", x"5b", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"40", x"5d", x"ff", x"fd", 
x"08", x"42", x"ff", x"ff", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"07", x"63", x"10", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"80", x"00", x"77", 
x"40", x"bd", x"ff", x"fb", 
x"47", x"a2", x"ff", x"fa", 
x"08", x"43", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f9", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"23", x"70", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"07", 
x"40", x"5d", x"ff", x"fa", 
x"08", x"42", x"ff", x"ff", 
x"40", x"7d", x"ff", x"ff", 
x"0a", x"03", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"40", x"90", x"00", x"05", 
x"40", x"b0", x"00", x"04", 
x"40", x"d0", x"00", x"03", 
x"40", x"f0", x"00", x"02", 
x"41", x"10", x"00", x"01", 
x"14", x"42", x"00", x"02", 
x"09", x"20", x"00", x"00", 
x"07", x"65", x"48", x"00", 
x"41", x"3b", x"00", x"00", 
x"09", x"40", x"00", x"37", 
x"c0", x"4a", x"00", x"00", 
x"40", x"63", x"00", x"07", 
x"09", x"40", x"00", x"00", 
x"07", x"63", x"50", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"08", x"60", x"00", x"00", 
x"07", x"67", x"18", x"00", 
x"c0", x"7b", x"00", x"00", 
x"98", x"63", x"00", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"67", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"98", x"84", x"00", x"00", 
x"08", x"60", x"00", x"02", 
x"07", x"67", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"98", x"a5", x"00", x"00", 
x"08", x"62", x"00", x"01", 
x"09", x"40", x"00", x"00", 
x"07", x"67", x"50", x"00", 
x"c0", x"db", x"00", x"00", 
x"09", x"40", x"00", x"03", 
x"09", x"60", x"00", x"38", 
x"c0", x"eb", x"00", x"00", 
x"47", x"a5", x"ff", x"ff", 
x"c7", x"a3", x"ff", x"fe", 
x"47", x"a7", x"ff", x"fd", 
x"47", x"a2", x"ff", x"fc", 
x"47", x"a9", x"ff", x"fb", 
x"47", x"a4", x"ff", x"fa", 
x"47", x"a3", x"ff", x"f9", 
x"c7", x"a2", x"ff", x"f8", 
x"47", x"a8", x"ff", x"f7", 
x"c7", x"a5", x"ff", x"f6", 
x"c7", x"a4", x"ff", x"f5", 
x"c7", x"a6", x"ff", x"f4", 
x"47", x"a6", x"ff", x"f3", 
x"08", x"4a", x"00", x"00", 
x"80", x"47", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"f2", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"f2", 
x"44", x"62", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"c0", x"5d", x"ff", x"f4", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"c0", x"5d", x"ff", x"f5", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"c0", x"7d", x"ff", x"f6", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"bd", x"ff", x"f7", 
x"47", x"a3", x"ff", x"f1", 
x"0a", x"05", x"00", x"00", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"23", x"db", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"c0", x"5d", x"ff", x"f8", 
x"c4", x"42", x"00", x"02", 
x"40", x"7d", x"ff", x"f1", 
x"44", x"43", x"00", x"01", 
x"40", x"7d", x"ff", x"f9", 
x"44", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"fb", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"43", x"00", x"01", 
x"40", x"bd", x"ff", x"fc", 
x"08", x"c5", x"00", x"02", 
x"08", x"e0", x"00", x"01", 
x"41", x"1d", x"ff", x"fd", 
x"07", x"68", x"38", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"e0", x"00", x"03", 
x"09", x"20", x"00", x"38", 
x"c0", x"89", x"00", x"00", 
x"47", x"a2", x"ff", x"f0", 
x"47", x"a6", x"ff", x"ef", 
x"c7", x"a3", x"ff", x"ee", 
x"08", x"47", x"00", x"00", 
x"80", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"ed", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"13", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"ed", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"ed", 
x"44", x"62", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"c0", x"5d", x"ff", x"fe", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"c0", x"7d", x"ff", x"ee", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"c0", x"7d", x"ff", x"f6", 
x"07", x"62", x"20", x"00", 
x"c7", x"63", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"bd", x"ff", x"f7", 
x"47", x"a3", x"ff", x"ec", 
x"0a", x"05", x"00", x"00", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"24", x"29", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"c0", x"5d", x"ff", x"f8", 
x"c4", x"42", x"00", x"02", 
x"40", x"7d", x"ff", x"ec", 
x"44", x"43", x"00", x"01", 
x"40", x"7d", x"ff", x"ef", 
x"44", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"f0", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"fb", 
x"08", x"62", x"00", x"02", 
x"40", x"bd", x"ff", x"fc", 
x"08", x"a5", x"00", x"03", 
x"08", x"c0", x"00", x"02", 
x"40", x"fd", x"ff", x"fd", 
x"07", x"67", x"30", x"00", 
x"c0", x"7b", x"00", x"00", 
x"08", x"c0", x"00", x"03", 
x"08", x"e0", x"00", x"38", 
x"c0", x"87", x"00", x"00", 
x"47", x"a3", x"ff", x"eb", 
x"47", x"a5", x"ff", x"ea", 
x"c7", x"a3", x"ff", x"e9", 
x"08", x"46", x"00", x"00", 
x"80", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"e8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"18", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"e8", 
x"0b", x"bd", x"ff", x"e7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"19", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"e8", 
x"44", x"62", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"c0", x"5d", x"ff", x"fe", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"c0", x"5d", x"ff", x"f5", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"c0", x"5d", x"ff", x"e9", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f3", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"f7", 
x"47", x"a3", x"ff", x"e7", 
x"0a", x"04", x"00", x"00", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"e6", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"24", x"78", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1a", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"c0", x"5d", x"ff", x"f8", 
x"c4", x"42", x"00", x"02", 
x"40", x"7d", x"ff", x"e7", 
x"44", x"43", x"00", x"01", 
x"40", x"7d", x"ff", x"ea", 
x"44", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"eb", 
x"40", x"9d", x"ff", x"fa", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fb", 
x"08", x"63", x"00", x"03", 
x"40", x"9d", x"ff", x"ff", 
x"07", x"64", x"10", x"00", 
x"47", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"05", 
x"40", x"b0", x"00", x"04", 
x"40", x"d0", x"00", x"03", 
x"40", x"f0", x"00", x"02", 
x"41", x"10", x"00", x"01", 
x"14", x"42", x"00", x"02", 
x"08", x"42", x"00", x"01", 
x"09", x"20", x"00", x"00", 
x"07", x"65", x"48", x"00", 
x"41", x"3b", x"00", x"00", 
x"09", x"40", x"00", x"37", 
x"c0", x"4a", x"00", x"00", 
x"41", x"43", x"00", x"07", 
x"09", x"60", x"00", x"00", 
x"07", x"6a", x"58", x"00", 
x"c0", x"7b", x"00", x"00", 
x"88", x"42", x"18", x"00", 
x"41", x"43", x"00", x"04", 
x"47", x"a5", x"ff", x"ff", 
x"47", x"a9", x"ff", x"fe", 
x"47", x"a4", x"ff", x"fd", 
x"47", x"a2", x"ff", x"fc", 
x"c7", x"a2", x"ff", x"fb", 
x"47", x"a8", x"ff", x"fa", 
x"47", x"a6", x"ff", x"f9", 
x"47", x"a7", x"ff", x"f8", 
x"47", x"a3", x"ff", x"f7", 
x"08", x"6a", x"00", x"00", 
x"08", x"47", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"79", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"40", x"00", x"32", 
x"c0", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f7", 
x"40", x"62", x"00", x"04", 
x"08", x"80", x"00", x"00", 
x"07", x"63", x"20", x"00", 
x"c0", x"9b", x"00", x"00", 
x"8c", x"63", x"20", x"00", 
x"8c", x"63", x"10", x"00", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f8", 
x"07", x"64", x"18", x"00", 
x"c0", x"9b", x"00", x"00", 
x"88", x"63", x"20", x"00", 
x"08", x"60", x"00", x"32", 
x"c0", x"83", x"00", x"00", 
x"40", x"62", x"00", x"04", 
x"08", x"a0", x"00", x"01", 
x"07", x"63", x"28", x"00", 
x"c0", x"bb", x"00", x"00", 
x"8c", x"84", x"28", x"00", 
x"8c", x"84", x"10", x"00", 
x"08", x"60", x"00", x"01", 
x"07", x"64", x"18", x"00", 
x"c0", x"bb", x"00", x"00", 
x"88", x"84", x"28", x"00", 
x"08", x"60", x"00", x"32", 
x"c0", x"a3", x"00", x"00", 
x"40", x"42", x"00", x"04", 
x"08", x"60", x"00", x"02", 
x"07", x"62", x"18", x"00", 
x"c0", x"db", x"00", x"00", 
x"8c", x"a5", x"30", x"00", 
x"8c", x"a5", x"10", x"00", 
x"08", x"40", x"00", x"02", 
x"07", x"64", x"10", x"00", 
x"c0", x"5b", x"00", x"00", 
x"88", x"a5", x"10", x"00", 
x"08", x"40", x"00", x"03", 
x"08", x"60", x"00", x"38", 
x"c0", x"43", x"00", x"00", 
x"c7", x"a5", x"ff", x"f6", 
x"c7", x"a4", x"ff", x"f5", 
x"c7", x"a3", x"ff", x"f4", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"a3", x"ff", x"f3", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"f3", 
x"44", x"62", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"c0", x"5d", x"ff", x"f4", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"01", 
x"c0", x"5d", x"ff", x"f5", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"80", x"00", x"02", 
x"c0", x"5d", x"ff", x"f6", 
x"07", x"62", x"20", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"40", x"9d", x"ff", x"f9", 
x"07", x"64", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fa", 
x"47", x"a3", x"ff", x"f2", 
x"0a", x"04", x"00", x"00", 
x"0b", x"63", x"00", x"00", 
x"08", x"62", x"00", x"00", 
x"08", x"5b", x"00", x"00", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"25", x"0c", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"c0", x"5d", x"ff", x"fb", 
x"c4", x"42", x"00", x"02", 
x"40", x"7d", x"ff", x"f2", 
x"44", x"43", x"00", x"01", 
x"40", x"7d", x"ff", x"fc", 
x"44", x"43", x"00", x"00", 
x"40", x"7d", x"ff", x"fe", 
x"40", x"9d", x"ff", x"fd", 
x"07", x"64", x"18", x"00", 
x"47", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"08", x"63", x"00", x"01", 
x"40", x"9d", x"ff", x"ff", 
x"07", x"64", x"10", x"00", 
x"47", x"63", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"70", x"00", x"03", 
x"40", x"90", x"00", x"02", 
x"40", x"b0", x"00", x"01", 
x"0b", x"60", x"00", x"00", 
x"2f", x"62", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"07", x"65", x"10", x"00", 
x"40", x"bb", x"00", x"00", 
x"40", x"c5", x"00", x"02", 
x"0b", x"60", x"00", x"02", 
x"20", x"db", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"40", x"c5", x"00", x"07", 
x"08", x"e0", x"00", x"00", 
x"07", x"66", x"38", x"00", 
x"c0", x"5b", x"00", x"00", 
x"08", x"c0", x"00", x"37", 
x"c0", x"66", x"00", x"00", 
x"ac", x"62", x"00", x"0e", 
x"40", x"c5", x"00", x"01", 
x"0b", x"60", x"00", x"01", 
x"20", x"db", x"00", x"07", 
x"0b", x"60", x"00", x"02", 
x"20", x"db", x"00", x"01", 
x"33", x"e0", x"00", x"00", 
x"0a", x"03", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"0a", x"04", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"40", x"90", x"00", x"10", 
x"40", x"b0", x"00", x"0f", 
x"40", x"d0", x"00", x"0e", 
x"40", x"f0", x"00", x"0d", 
x"41", x"10", x"00", x"0c", 
x"41", x"30", x"00", x"0b", 
x"41", x"50", x"00", x"0a", 
x"41", x"70", x"00", x"09", 
x"41", x"90", x"00", x"08", 
x"41", x"b0", x"00", x"07", 
x"41", x"d0", x"00", x"06", 
x"41", x"f0", x"00", x"05", 
x"47", x"a8", x"ff", x"ff", 
x"41", x"10", x"00", x"04", 
x"47", x"aa", x"ff", x"fe", 
x"41", x"50", x"00", x"03", 
x"47", x"a6", x"ff", x"fd", 
x"40", x"d0", x"00", x"02", 
x"47", x"ac", x"ff", x"fc", 
x"41", x"90", x"00", x"01", 
x"47", x"ae", x"ff", x"fb", 
x"09", x"c0", x"00", x"00", 
x"07", x"68", x"70", x"00", 
x"47", x"62", x"00", x"00", 
x"09", x"c0", x"00", x"01", 
x"07", x"68", x"70", x"00", 
x"47", x"63", x"00", x"00", 
x"09", x"c0", x"00", x"00", 
x"47", x"ab", x"ff", x"fa", 
x"19", x"62", x"00", x"01", 
x"07", x"6a", x"70", x"00", 
x"47", x"6b", x"00", x"00", 
x"09", x"60", x"00", x"01", 
x"18", x"63", x"00", x"01", 
x"07", x"6a", x"58", x"00", 
x"47", x"63", x"00", x"00", 
x"08", x"60", x"00", x"00", 
x"09", x"40", x"00", x"19", 
x"c0", x"4a", x"00", x"00", 
x"b4", x"62", x"00", x"00", 
x"93", x"63", x"00", x"00", 
x"8c", x"42", x"d8", x"00", 
x"07", x"67", x"18", x"00", 
x"c7", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"07", x"68", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"47", x"ad", x"ff", x"f9", 
x"47", x"a5", x"ff", x"f8", 
x"47", x"af", x"ff", x"f7", 
x"47", x"ac", x"ff", x"f6", 
x"47", x"a6", x"ff", x"f5", 
x"47", x"a4", x"ff", x"f4", 
x"47", x"a9", x"ff", x"f3", 
x"47", x"a8", x"ff", x"f2", 
x"47", x"a2", x"ff", x"f1", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"92", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"08", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f1", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f2", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"63", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"e3", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f2", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"47", x"a2", x"ff", x"f0", 
x"47", x"a3", x"ff", x"ef", 
x"0b", x"bd", x"ff", x"ee", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"92", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"12", 
x"08", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"ef", 
x"0b", x"bd", x"ff", x"ee", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"12", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f2", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"63", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"ee", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"e3", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"12", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f2", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"47", x"a2", x"ff", x"ee", 
x"47", x"a3", x"ff", x"ed", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"92", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"08", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"ed", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"08", x"60", x"00", x"00", 
x"40", x"9d", x"ff", x"f2", 
x"07", x"64", x"18", x"00", 
x"40", x"7b", x"00", x"00", 
x"08", x"63", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"20", x"e3", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"40", x"7d", x"ff", x"f3", 
x"47", x"a2", x"ff", x"ec", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"25", x"d0", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"40", x"5d", x"ff", x"f4", 
x"0a", x"02", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"25", x"d9", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f5", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"25", x"e3", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"40", x"00", x"09", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"bd", x"ff", x"f6", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"25", x"ef", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"40", x"00", x"04", 
x"40", x"7d", x"ff", x"f7", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"25", x"f9", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"40", x"5d", x"ff", x"f8", 
x"40", x"7d", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"00", x"03", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"9d", x"ff", x"fc", 
x"40", x"bd", x"ff", x"fb", 
x"08", x"62", x"00", x"00", 
x"0a", x"05", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"26", x"11", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"40", x"00", x"00", 
x"40", x"7d", x"ff", x"fa", 
x"07", x"63", x"10", x"00", 
x"40", x"5b", x"00", x"00", 
x"08", x"42", x"ff", x"ff", 
x"40", x"7d", x"ff", x"fd", 
x"0a", x"03", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"26", x"1f", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"40", x"5d", x"ff", x"ee", 
x"40", x"bd", x"ff", x"fe", 
x"0a", x"05", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"26", x"2b", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"40", x"00", x"00", 
x"08", x"c0", x"00", x"02", 
x"40", x"7d", x"ff", x"f0", 
x"40", x"9d", x"ff", x"ee", 
x"40", x"bd", x"ff", x"ec", 
x"40", x"fd", x"ff", x"ff", 
x"0a", x"07", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"33", x"60", x"00", x"00", 
x"0b", x"a0", x"03", x"ff", 
x"17", x"bd", x"00", x"0a", 
x"0b", x"bd", x"03", x"ff", 
x"0b", x"80", x"03", x"ff", 
x"08", x"40", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"60", x"00", x"3c", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"00", 
x"08", x"c0", x"00", x"00", 
x"08", x"e0", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"09", x"3c", x"00", x"00", 
x"0b", x"9c", x"00", x"0b", 
x"45", x"22", x"00", x"0a", 
x"45", x"22", x"00", x"09", 
x"45", x"22", x"00", x"08", 
x"45", x"22", x"00", x"07", 
x"45", x"28", x"00", x"06", 
x"45", x"22", x"00", x"05", 
x"45", x"22", x"00", x"04", 
x"45", x"27", x"00", x"03", 
x"45", x"26", x"00", x"02", 
x"45", x"25", x"00", x"01", 
x"45", x"24", x"00", x"00", 
x"08", x"43", x"00", x"00", 
x"08", x"69", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"fe", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"fd", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"fc", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"26", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"fb", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"fa", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"06", 
x"08", x"60", x"00", x"32", 
x"08", x"80", x"00", x"01", 
x"08", x"a0", x"ff", x"ff", 
x"47", x"a2", x"ff", x"fa", 
x"47", x"a3", x"ff", x"f9", 
x"08", x"65", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"08", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f9", 
x"0b", x"bd", x"ff", x"f8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"08", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"01", 
x"08", x"a0", x"00", x"00", 
x"07", x"62", x"28", x"00", 
x"40", x"bb", x"00", x"00", 
x"47", x"a2", x"ff", x"f8", 
x"47", x"a3", x"ff", x"f7", 
x"08", x"65", x"00", x"00", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"62", x"00", x"00", 
x"40", x"5d", x"ff", x"f7", 
x"0b", x"bd", x"ff", x"f6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0a", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"f6", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0b", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"f5", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0c", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"2d", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"f4", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0d", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"f3", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0e", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"f2", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"f1", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"0f", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"f1", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"f0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"10", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"f0", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"ef", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"11", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"ef", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"ee", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"12", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"ee", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"ed", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"13", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"ed", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"ec", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"14", 
x"08", x"60", x"00", x"02", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"ec", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"eb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"15", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"eb", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"ea", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"16", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"ea", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e9", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"17", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e9", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e8", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"18", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e8", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e7", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"19", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e7", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e6", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1a", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e6", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e5", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1b", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e5", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e4", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1c", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e4", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e3", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1d", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"47", x"a3", x"ff", x"e3", 
x"0b", x"bd", x"ff", x"e2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1e", 
x"08", x"60", x"00", x"00", 
x"08", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"82", x"00", x"01", 
x"40", x"5d", x"ff", x"e3", 
x"44", x"82", x"00", x"00", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"e2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1e", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"05", 
x"0b", x"bd", x"ff", x"e2", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1e", 
x"08", x"60", x"00", x"00", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e2", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e1", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"1f", 
x"08", x"60", x"00", x"03", 
x"08", x"80", x"00", x"38", 
x"c0", x"44", x"00", x"00", 
x"47", x"a2", x"ff", x"e1", 
x"08", x"43", x"00", x"00", 
x"0b", x"bd", x"ff", x"e0", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"20", 
x"08", x"60", x"00", x"3c", 
x"40", x"9d", x"ff", x"e1", 
x"47", x"a2", x"ff", x"e0", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"df", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"21", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"e0", 
x"44", x"62", x"00", x"00", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"47", x"a3", x"ff", x"df", 
x"08", x"44", x"00", x"00", 
x"0b", x"bd", x"ff", x"de", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"37", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"22", 
x"08", x"62", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"47", x"a3", x"ff", x"de", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"44", x"62", x"00", x"01", 
x"40", x"5d", x"ff", x"de", 
x"44", x"62", x"00", x"00", 
x"08", x"40", x"00", x"b4", 
x"08", x"80", x"00", x"00", 
x"08", x"a0", x"00", x"38", 
x"c0", x"45", x"00", x"00", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"c4", x"a2", x"00", x"02", 
x"44", x"a3", x"00", x"01", 
x"44", x"a4", x"00", x"00", 
x"08", x"65", x"00", x"00", 
x"0b", x"bd", x"ff", x"dd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"23", 
x"08", x"60", x"00", x"01", 
x"08", x"80", x"00", x"00", 
x"47", x"a2", x"ff", x"dd", 
x"08", x"43", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"dc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"2f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"24", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"06", 
x"08", x"80", x"01", x"22", 
x"44", x"64", x"00", x"00", 
x"40", x"9d", x"ff", x"fc", 
x"44", x"64", x"00", x"05", 
x"40", x"bd", x"ff", x"e5", 
x"44", x"65", x"00", x"04", 
x"40", x"dd", x"ff", x"e6", 
x"44", x"66", x"00", x"03", 
x"40", x"fd", x"ff", x"e7", 
x"44", x"67", x"00", x"02", 
x"41", x"1d", x"ff", x"fd", 
x"44", x"68", x"00", x"01", 
x"09", x"1c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"20", x"01", x"cf", 
x"45", x"09", x"00", x"00", 
x"41", x"3d", x"ff", x"fb", 
x"45", x"09", x"00", x"02", 
x"41", x"5d", x"ff", x"fa", 
x"45", x"0a", x"00", x"01", 
x"09", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"80", x"02", x"d3", 
x"45", x"6c", x"00", x"00", 
x"41", x"9d", x"ff", x"fe", 
x"45", x"6c", x"00", x"01", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"c0", x"05", x"31", 
x"45", x"ae", x"00", x"00", 
x"45", x"ab", x"00", x"02", 
x"41", x"7d", x"ff", x"ff", 
x"45", x"ab", x"00", x"01", 
x"09", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"e0", x"05", x"9e", 
x"45", x"cf", x"00", x"00", 
x"41", x"fd", x"ff", x"f8", 
x"45", x"cf", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"07", 
x"08", x"a0", x"05", x"ca", 
x"44", x"c5", x"00", x"00", 
x"44", x"c3", x"00", x"06", 
x"44", x"cd", x"00", x"05", 
x"44", x"c8", x"00", x"04", 
x"44", x"ce", x"00", x"03", 
x"40", x"7d", x"ff", x"f6", 
x"44", x"c3", x"00", x"02", 
x"44", x"cf", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"00", x"06", x"28", 
x"44", x"a8", x"00", x"00", 
x"41", x"1d", x"ff", x"f5", 
x"44", x"a8", x"00", x"01", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"c0", x"06", x"c3", 
x"45", x"ae", x"00", x"00", 
x"45", x"a5", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"c0", x"07", x"6a", 
x"44", x"ae", x"00", x"00", 
x"44", x"a8", x"00", x"01", 
x"09", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"05", 
x"47", x"a6", x"ff", x"dc", 
x"08", x"c0", x"07", x"f9", 
x"45", x"c6", x"00", x"00", 
x"45", x"c5", x"00", x"04", 
x"45", x"cd", x"00", x"03", 
x"45", x"c8", x"00", x"02", 
x"45", x"cc", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"c0", x"08", x"4f", 
x"44", x"a6", x"00", x"00", 
x"44", x"a8", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"a0", x"08", x"e9", 
x"44", x"cd", x"00", x"00", 
x"44", x"c8", x"00", x"01", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"e0", x"09", x"05", 
x"45", x"a7", x"00", x"00", 
x"45", x"a8", x"00", x"01", 
x"08", x"fc", x"00", x"00", 
x"0b", x"9c", x"00", x"05", 
x"08", x"80", x"09", x"7d", 
x"44", x"e4", x"00", x"00", 
x"44", x"e6", x"00", x"04", 
x"44", x"ed", x"00", x"03", 
x"44", x"e5", x"00", x"02", 
x"44", x"ec", x"00", x"01", 
x"08", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"c0", x"09", x"b2", 
x"44", x"86", x"00", x"00", 
x"44", x"88", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"a0", x"09", x"c7", 
x"44", x"cd", x"00", x"00", 
x"44", x"c8", x"00", x"01", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"05", 
x"09", x"40", x"0a", x"05", 
x"45", x"aa", x"00", x"00", 
x"45", x"a4", x"00", x"04", 
x"45", x"a6", x"00", x"03", 
x"45", x"a5", x"00", x"02", 
x"45", x"ac", x"00", x"01", 
x"08", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"a0", x"0c", x"63", 
x"44", x"85", x"00", x"00", 
x"44", x"8c", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"c0", x"0c", x"af", 
x"44", x"a6", x"00", x"00", 
x"44", x"ac", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"40", x"0d", x"ab", 
x"44", x"ca", x"00", x"00", 
x"44", x"cc", x"00", x"01", 
x"09", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"08", 
x"47", x"a4", x"ff", x"db", 
x"08", x"80", x"0d", x"e7", 
x"45", x"44", x"00", x"00", 
x"45", x"47", x"00", x"07", 
x"45", x"48", x"00", x"06", 
x"45", x"4c", x"00", x"05", 
x"40", x"9d", x"ff", x"df", 
x"45", x"44", x"00", x"04", 
x"45", x"49", x"00", x"03", 
x"41", x"3d", x"ff", x"f2", 
x"45", x"49", x"00", x"02", 
x"45", x"46", x"00", x"01", 
x"09", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"47", x"a2", x"ff", x"da", 
x"08", x"40", x"0e", x"7a", 
x"45", x"62", x"00", x"00", 
x"45", x"6a", x"00", x"02", 
x"45", x"6f", x"00", x"01", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"06", 
x"09", x"40", x"0e", x"9c", 
x"44", x"4a", x"00", x"00", 
x"44", x"47", x"00", x"05", 
x"44", x"48", x"00", x"04", 
x"44", x"4b", x"00", x"03", 
x"44", x"44", x"00", x"02", 
x"44", x"49", x"00", x"01", 
x"08", x"fc", x"00", x"00", 
x"0b", x"9c", x"00", x"0a", 
x"09", x"40", x"0f", x"13", 
x"44", x"ea", x"00", x"00", 
x"41", x"5d", x"ff", x"f3", 
x"44", x"ea", x"00", x"09", 
x"41", x"7d", x"ff", x"e9", 
x"44", x"eb", x"00", x"08", 
x"44", x"e8", x"00", x"07", 
x"44", x"ee", x"00", x"06", 
x"44", x"ec", x"00", x"05", 
x"40", x"9d", x"ff", x"f4", 
x"44", x"e4", x"00", x"04", 
x"44", x"e9", x"00", x"03", 
x"47", x"a5", x"ff", x"d9", 
x"40", x"bd", x"ff", x"f1", 
x"44", x"e5", x"00", x"02", 
x"44", x"e6", x"00", x"01", 
x"47", x"a2", x"ff", x"d8", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"47", x"a6", x"ff", x"d7", 
x"08", x"c0", x"10", x"03", 
x"44", x"46", x"00", x"00", 
x"44", x"47", x"00", x"02", 
x"44", x"4f", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"08", 
x"08", x"a0", x"10", x"3f", 
x"44", x"c5", x"00", x"00", 
x"44", x"ca", x"00", x"07", 
x"44", x"cb", x"00", x"06", 
x"44", x"c8", x"00", x"05", 
x"44", x"ce", x"00", x"04", 
x"44", x"c2", x"00", x"03", 
x"44", x"c7", x"00", x"02", 
x"44", x"cf", x"00", x"01", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"04", 
x"08", x"a0", x"10", x"e1", 
x"44", x"45", x"00", x"00", 
x"44", x"46", x"00", x"03", 
x"44", x"4a", x"00", x"02", 
x"44", x"43", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"0a", 
x"08", x"c0", x"11", x"09", 
x"44", x"a6", x"00", x"00", 
x"44", x"aa", x"00", x"09", 
x"40", x"dd", x"ff", x"e8", 
x"44", x"a6", x"00", x"08", 
x"44", x"ad", x"00", x"07", 
x"44", x"a8", x"00", x"06", 
x"44", x"ac", x"00", x"05", 
x"44", x"a4", x"00", x"04", 
x"44", x"a9", x"00", x"03", 
x"40", x"fd", x"ff", x"f1", 
x"44", x"a7", x"00", x"02", 
x"41", x"dd", x"ff", x"d7", 
x"44", x"ae", x"00", x"01", 
x"09", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"47", x"a2", x"ff", x"d6", 
x"08", x"40", x"11", x"fa", 
x"45", x"c2", x"00", x"00", 
x"45", x"c5", x"00", x"02", 
x"45", x"cf", x"00", x"01", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"07", 
x"09", x"80", x"12", x"36", 
x"44", x"4c", x"00", x"00", 
x"44", x"4a", x"00", x"06", 
x"44", x"4d", x"00", x"05", 
x"44", x"48", x"00", x"04", 
x"44", x"4e", x"00", x"03", 
x"44", x"45", x"00", x"02", 
x"44", x"4f", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"04", 
x"09", x"00", x"12", x"d6", 
x"44", x"a8", x"00", x"00", 
x"44", x"a2", x"00", x"03", 
x"44", x"aa", x"00", x"02", 
x"44", x"a3", x"00", x"01", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"00", x"12", x"fe", 
x"44", x"48", x"00", x"00", 
x"41", x"1d", x"ff", x"f0", 
x"44", x"48", x"00", x"02", 
x"44", x"44", x"00", x"01", 
x"09", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"a0", x"13", x"27", 
x"45", x"8d", x"00", x"00", 
x"45", x"88", x"00", x"01", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"c0", x"13", x"41", 
x"45", x"ae", x"00", x"00", 
x"45", x"a8", x"00", x"02", 
x"45", x"a9", x"00", x"01", 
x"09", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"e0", x"13", x"b5", 
x"45", x"cf", x"00", x"00", 
x"41", x"fd", x"ff", x"ef", 
x"45", x"cf", x"00", x"01", 
x"47", x"ac", x"ff", x"d5", 
x"09", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"47", x"a2", x"ff", x"d4", 
x"08", x"40", x"15", x"2d", 
x"45", x"82", x"00", x"00", 
x"45", x"8f", x"00", x"02", 
x"40", x"5d", x"ff", x"ed", 
x"45", x"82", x"00", x"01", 
x"47", x"ad", x"ff", x"d3", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"09", 
x"09", x"20", x"15", x"7b", 
x"45", x"a9", x"00", x"00", 
x"41", x"3d", x"ff", x"d8", 
x"45", x"a9", x"00", x"08", 
x"40", x"5d", x"ff", x"dd", 
x"45", x"a2", x"00", x"07", 
x"45", x"a3", x"00", x"06", 
x"45", x"a8", x"00", x"05", 
x"45", x"a5", x"00", x"04", 
x"45", x"a4", x"00", x"03", 
x"45", x"a7", x"00", x"02", 
x"45", x"ac", x"00", x"01", 
x"08", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"19", 
x"47", x"a5", x"ff", x"d2", 
x"08", x"a0", x"16", x"06", 
x"44", x"45", x"00", x"00", 
x"44", x"4e", x"00", x"18", 
x"44", x"4d", x"00", x"17", 
x"44", x"4a", x"00", x"16", 
x"44", x"4f", x"00", x"15", 
x"44", x"46", x"00", x"14", 
x"44", x"4b", x"00", x"13", 
x"44", x"49", x"00", x"12", 
x"40", x"bd", x"ff", x"d9", 
x"44", x"45", x"00", x"11", 
x"41", x"5d", x"ff", x"ed", 
x"44", x"4a", x"00", x"10", 
x"44", x"43", x"00", x"0f", 
x"41", x"bd", x"ff", x"fe", 
x"44", x"4d", x"00", x"0e", 
x"44", x"48", x"00", x"0d", 
x"41", x"7d", x"ff", x"da", 
x"44", x"4b", x"00", x"0c", 
x"41", x"7d", x"ff", x"ff", 
x"44", x"4b", x"00", x"0b", 
x"41", x"5d", x"ff", x"fb", 
x"44", x"4a", x"00", x"0a", 
x"41", x"7d", x"ff", x"d6", 
x"44", x"4b", x"00", x"09", 
x"44", x"44", x"00", x"08", 
x"40", x"9d", x"ff", x"f2", 
x"44", x"44", x"00", x"07", 
x"44", x"47", x"00", x"06", 
x"41", x"7d", x"ff", x"d3", 
x"44", x"4b", x"00", x"05", 
x"40", x"bd", x"ff", x"d4", 
x"44", x"45", x"00", x"04", 
x"40", x"dd", x"ff", x"d5", 
x"44", x"46", x"00", x"03", 
x"40", x"dd", x"ff", x"fa", 
x"44", x"46", x"00", x"02", 
x"44", x"4c", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"0f", 
x"09", x"80", x"17", x"cf", 
x"44", x"cc", x"00", x"00", 
x"44", x"ce", x"00", x"0e", 
x"44", x"cf", x"00", x"0d", 
x"44", x"c9", x"00", x"0c", 
x"44", x"c3", x"00", x"0b", 
x"44", x"cd", x"00", x"0a", 
x"44", x"c8", x"00", x"09", 
x"44", x"ca", x"00", x"08", 
x"40", x"7d", x"ff", x"d2", 
x"44", x"c3", x"00", x"07", 
x"44", x"c4", x"00", x"06", 
x"44", x"c7", x"00", x"05", 
x"44", x"cb", x"00", x"04", 
x"44", x"c5", x"00", x"03", 
x"40", x"7d", x"ff", x"d5", 
x"44", x"c3", x"00", x"02", 
x"40", x"7d", x"ff", x"ee", 
x"44", x"c3", x"00", x"01", 
x"08", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"a0", x"18", x"dd", 
x"44", x"85", x"00", x"00", 
x"44", x"86", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"06", 
x"08", x"c0", x"19", x"2a", 
x"44", x"a6", x"00", x"00", 
x"40", x"dd", x"ff", x"e8", 
x"44", x"a6", x"00", x"05", 
x"40", x"fd", x"ff", x"d9", 
x"44", x"a7", x"00", x"04", 
x"41", x"1d", x"ff", x"ff", 
x"44", x"a8", x"00", x"03", 
x"44", x"a4", x"00", x"02", 
x"41", x"3d", x"ff", x"e2", 
x"44", x"a9", x"00", x"01", 
x"09", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"04", 
x"09", x"80", x"1b", x"ec", 
x"45", x"6c", x"00", x"00", 
x"45", x"65", x"00", x"03", 
x"40", x"bd", x"ff", x"ed", 
x"45", x"65", x"00", x"02", 
x"45", x"63", x"00", x"01", 
x"09", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"c0", x"1c", x"22", 
x"45", x"8e", x"00", x"00", 
x"45", x"85", x"00", x"02", 
x"45", x"83", x"00", x"01", 
x"09", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"e0", x"1c", x"7d", 
x"45", x"cf", x"00", x"00", 
x"45", x"cb", x"00", x"01", 
x"09", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"e0", x"1c", x"a0", 
x"45", x"6f", x"00", x"00", 
x"41", x"fd", x"ff", x"ec", 
x"45", x"6f", x"00", x"01", 
x"09", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"40", x"1c", x"e2", 
x"45", x"aa", x"00", x"00", 
x"45", x"ae", x"00", x"02", 
x"45", x"ac", x"00", x"01", 
x"09", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"80", x"1d", x"34", 
x"45", x"4c", x"00", x"00", 
x"45", x"4f", x"00", x"01", 
x"09", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"47", x"aa", x"ff", x"d1", 
x"09", x"40", x"1d", x"6f", 
x"45", x"8a", x"00", x"00", 
x"45", x"85", x"00", x"01", 
x"09", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"07", 
x"47", x"ae", x"ff", x"d0", 
x"09", x"c0", x"1e", x"21", 
x"45", x"4e", x"00", x"00", 
x"45", x"46", x"00", x"06", 
x"45", x"47", x"00", x"05", 
x"45", x"48", x"00", x"04", 
x"45", x"44", x"00", x"03", 
x"45", x"49", x"00", x"02", 
x"45", x"43", x"00", x"01", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"0a", 
x"08", x"80", x"1e", x"8f", 
x"44", x"64", x"00", x"00", 
x"40", x"9d", x"ff", x"fc", 
x"44", x"64", x"00", x"09", 
x"44", x"62", x"00", x"08", 
x"40", x"5d", x"ff", x"e9", 
x"44", x"62", x"00", x"07", 
x"40", x"5d", x"ff", x"e7", 
x"44", x"62", x"00", x"06", 
x"40", x"5d", x"ff", x"ea", 
x"44", x"62", x"00", x"05", 
x"44", x"65", x"00", x"04", 
x"40", x"9d", x"ff", x"e4", 
x"44", x"64", x"00", x"03", 
x"44", x"6a", x"00", x"02", 
x"40", x"9d", x"ff", x"eb", 
x"44", x"64", x"00", x"01", 
x"08", x"dc", x"00", x"00", 
x"0b", x"9c", x"00", x"07", 
x"08", x"e0", x"1f", x"35", 
x"44", x"c7", x"00", x"00", 
x"40", x"fd", x"ff", x"e5", 
x"44", x"c7", x"00", x"06", 
x"40", x"fd", x"ff", x"e6", 
x"44", x"c7", x"00", x"05", 
x"44", x"c2", x"00", x"04", 
x"44", x"c3", x"00", x"03", 
x"44", x"cf", x"00", x"02", 
x"44", x"c4", x"00", x"01", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"07", 
x"08", x"e0", x"1f", x"67", 
x"44", x"67", x"00", x"00", 
x"44", x"6c", x"00", x"06", 
x"44", x"6d", x"00", x"05", 
x"44", x"65", x"00", x"04", 
x"44", x"6b", x"00", x"03", 
x"44", x"6f", x"00", x"02", 
x"40", x"bd", x"ff", x"d0", 
x"44", x"65", x"00", x"01", 
x"08", x"bc", x"00", x"00", 
x"0b", x"9c", x"00", x"04", 
x"08", x"e0", x"1f", x"d8", 
x"44", x"a7", x"00", x"00", 
x"44", x"a3", x"00", x"03", 
x"44", x"a6", x"00", x"02", 
x"44", x"af", x"00", x"01", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"08", x"e0", x"21", x"03", 
x"44", x"67", x"00", x"00", 
x"44", x"69", x"00", x"01", 
x"08", x"fc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"40", x"21", x"cb", 
x"44", x"ea", x"00", x"00", 
x"44", x"e3", x"00", x"01", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"40", x"22", x"1e", 
x"44", x"6a", x"00", x"00", 
x"44", x"67", x"00", x"01", 
x"08", x"fc", x"00", x"00", 
x"0b", x"9c", x"00", x"02", 
x"09", x"40", x"22", x"4a", 
x"44", x"ea", x"00", x"00", 
x"44", x"e8", x"00", x"01", 
x"09", x"5c", x"00", x"00", 
x"0b", x"9c", x"00", x"04", 
x"09", x"60", x"22", x"97", 
x"45", x"4b", x"00", x"00", 
x"45", x"48", x"00", x"03", 
x"45", x"49", x"00", x"02", 
x"45", x"47", x"00", x"01", 
x"08", x"fc", x"00", x"00", 
x"0b", x"9c", x"00", x"03", 
x"09", x"60", x"22", x"fa", 
x"44", x"eb", x"00", x"00", 
x"44", x"e8", x"00", x"02", 
x"41", x"7d", x"ff", x"db", 
x"44", x"eb", x"00", x"01", 
x"09", x"9c", x"00", x"00", 
x"0b", x"9c", x"00", x"05", 
x"09", x"a0", x"23", x"34", 
x"45", x"8d", x"00", x"00", 
x"45", x"88", x"00", x"04", 
x"45", x"8b", x"00", x"03", 
x"45", x"87", x"00", x"02", 
x"45", x"89", x"00", x"01", 
x"08", x"fc", x"00", x"00", 
x"0b", x"9c", x"00", x"06", 
x"09", x"20", x"23", x"78", 
x"44", x"e9", x"00", x"00", 
x"41", x"3d", x"ff", x"dd", 
x"44", x"e9", x"00", x"05", 
x"41", x"bd", x"ff", x"da", 
x"44", x"ed", x"00", x"04", 
x"44", x"e8", x"00", x"03", 
x"41", x"dd", x"ff", x"fb", 
x"44", x"ee", x"00", x"02", 
x"44", x"eb", x"00", x"01", 
x"47", x"a3", x"ff", x"cf", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"06", 
x"47", x"aa", x"ff", x"ce", 
x"09", x"40", x"24", x"8d", 
x"44", x"6a", x"00", x"00", 
x"44", x"69", x"00", x"05", 
x"44", x"6d", x"00", x"04", 
x"44", x"68", x"00", x"03", 
x"44", x"6e", x"00", x"02", 
x"44", x"6b", x"00", x"01", 
x"09", x"3c", x"00", x"00", 
x"0b", x"9c", x"00", x"04", 
x"09", x"40", x"25", x"20", 
x"45", x"2a", x"00", x"00", 
x"45", x"23", x"00", x"03", 
x"45", x"27", x"00", x"02", 
x"40", x"7d", x"ff", x"fe", 
x"45", x"23", x"00", x"01", 
x"08", x"7c", x"00", x"00", 
x"0b", x"9c", x"00", x"11", 
x"08", x"e0", x"25", x"42", 
x"44", x"67", x"00", x"00", 
x"40", x"fd", x"ff", x"d1", 
x"44", x"67", x"00", x"10", 
x"40", x"fd", x"ff", x"e0", 
x"44", x"67", x"00", x"0f", 
x"44", x"69", x"00", x"0e", 
x"44", x"62", x"00", x"0d", 
x"44", x"65", x"00", x"0c", 
x"40", x"5d", x"ff", x"dc", 
x"44", x"62", x"00", x"0b", 
x"44", x"66", x"00", x"0a", 
x"44", x"68", x"00", x"09", 
x"40", x"5d", x"ff", x"df", 
x"44", x"62", x"00", x"08", 
x"44", x"6e", x"00", x"07", 
x"44", x"6b", x"00", x"06", 
x"44", x"6c", x"00", x"05", 
x"44", x"6f", x"00", x"04", 
x"44", x"64", x"00", x"03", 
x"40", x"5d", x"ff", x"ce", 
x"44", x"62", x"00", x"02", 
x"40", x"5d", x"ff", x"cf", 
x"44", x"62", x"00", x"01", 
x"08", x"40", x"00", x"80", 
x"08", x"80", x"00", x"80", 
x"0a", x"03", x"00", x"00", 
x"08", x"64", x"00", x"00", 
x"0b", x"bd", x"ff", x"cd", 
x"47", x"bf", x"00", x"00", 
x"43", x"70", x"00", x"00", 
x"0f", x"e0", x"2a", x"2b", 
x"33", x"60", x"00", x"00", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"33", 
x"08", x"40", x"00", x"00", 
x"7c", x"00", x"00", x"00", 
x"05", x"00", x"10", x"00", 
x"04", x"40", x"e0", x"00", 
x"21", x"00", x"00", x"04", 
x"47", x"83", x"00", x"00", 
x"09", x"08", x"ff", x"ff", 
x"0b", x"9c", x"00", x"01", 
x"20", x"00", x"ff", x"fb", 
x"33", x"e0", x"00", x"00", 
x"05", x"00", x"10", x"00", 
x"04", x"40", x"e0", x"00", 
x"21", x"00", x"00", x"04", 
x"c7", x"82", x"00", x"00", 
x"09", x"08", x"ff", x"ff", 
x"0b", x"9c", x"00", x"01", 
x"20", x"00", x"ff", x"fb", 
x"33", x"e0", x"00", x"00", 
x"05", x"00", x"10", x"00", 
x"14", x"48", x"ff", x"fe", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fd", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"ff", 
x"04", x"42", x"40", x"00", 
x"14", x"42", x"ff", x"fc", 
x"33", x"e0", x"00", x"00", 
x"09", x"00", x"00", x"0a", 
x"75", x"00", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"74", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"2c", x"02", x"00", x"03", 
x"09", x"00", x"00", x"2d", 
x"75", x"00", x"00", x"00", 
x"10", x"40", x"10", x"00", 
x"09", x"80", x"00", x"08", 
x"05", x"00", x"00", x"00", 
x"05", x"20", x"00", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"a8", x"ff", x"fe", 
x"47", x"a9", x"ff", x"fd", 
x"47", x"ac", x"ff", x"fc", 
x"0b", x"bd", x"ff", x"fb", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"3f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"05", 
x"41", x"1d", x"ff", x"ff", 
x"41", x"9d", x"ff", x"fc", 
x"15", x"42", x"00", x"01", 
x"15", x"62", x"00", x"03", 
x"05", x"4a", x"58", x"00", 
x"11", x"48", x"50", x"00", 
x"09", x"4a", x"00", x"30", 
x"41", x"1d", x"ff", x"fe", 
x"41", x"3d", x"ff", x"fd", 
x"15", x"29", x"00", x"08", 
x"15", x"68", x"ff", x"e8", 
x"05", x"29", x"58", x"00", 
x"15", x"08", x"00", x"08", 
x"05", x"08", x"50", x"00", 
x"20", x"40", x"00", x"17", 
x"09", x"8c", x"ff", x"ff", 
x"21", x"80", x"00", x"01", 
x"20", x"00", x"ff", x"e5", 
x"47", x"a2", x"ff", x"ff", 
x"47", x"a8", x"ff", x"fe", 
x"47", x"a9", x"ff", x"fd", 
x"0b", x"bd", x"ff", x"fc", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"3f", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"04", 
x"41", x"1d", x"ff", x"ff", 
x"15", x"42", x"00", x"01", 
x"15", x"62", x"00", x"03", 
x"05", x"4a", x"58", x"00", 
x"11", x"48", x"50", x"00", 
x"09", x"4a", x"00", x"30", 
x"20", x"40", x"00", x"02", 
x"08", x"42", x"00", x"30", 
x"74", x"40", x"00", x"00", 
x"75", x"40", x"00", x"00", 
x"41", x"1d", x"ff", x"fe", 
x"41", x"3d", x"ff", x"fd", 
x"75", x"00", x"00", x"00", 
x"15", x"08", x"ff", x"f8", 
x"21", x"00", x"00", x"12", 
x"75", x"00", x"00", x"00", 
x"15", x"08", x"ff", x"f8", 
x"21", x"00", x"00", x"0f", 
x"75", x"00", x"00", x"00", 
x"15", x"08", x"ff", x"f8", 
x"21", x"00", x"00", x"0c", 
x"75", x"00", x"00", x"00", 
x"21", x"20", x"00", x"0a", 
x"75", x"20", x"00", x"00", 
x"15", x"29", x"ff", x"f8", 
x"21", x"20", x"00", x"07", 
x"75", x"20", x"00", x"00", 
x"15", x"29", x"ff", x"f8", 
x"21", x"20", x"00", x"04", 
x"75", x"20", x"00", x"00", 
x"15", x"29", x"ff", x"f8", 
x"21", x"20", x"00", x"01", 
x"75", x"20", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"15", x"42", x"ff", x"e8", 
x"75", x"40", x"00", x"00", 
x"15", x"42", x"ff", x"f0", 
x"75", x"40", x"00", x"00", 
x"15", x"42", x"ff", x"f8", 
x"75", x"40", x"00", x"00", 
x"74", x"40", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"c7", x"a2", x"ff", x"ff", 
x"41", x"1d", x"ff", x"ff", 
x"15", x"48", x"ff", x"e8", 
x"75", x"40", x"00", x"00", 
x"15", x"48", x"ff", x"f0", 
x"75", x"40", x"00", x"00", 
x"15", x"48", x"ff", x"f8", 
x"75", x"40", x"00", x"00", 
x"75", x"00", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"09", x"20", x"00", x"30", 
x"09", x"40", x"00", x"39", 
x"08", x"60", x"00", x"00", 
x"09", x"60", x"00", x"2d", 
x"78", x"60", x"00", x"00", 
x"20", x"6b", x"00", x"04", 
x"2d", x"23", x"00", x"01", 
x"20", x"00", x"ff", x"fc", 
x"2c", x"6a", x"00", x"04", 
x"20", x"00", x"ff", x"fa", 
x"09", x"00", x"00", x"01", 
x"08", x"40", x"00", x"00", 
x"20", x"00", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"08", x"43", x"ff", x"d0", 
x"78", x"60", x"00", x"00", 
x"28", x"69", x"00", x"07", 
x"29", x"43", x"00", x"06", 
x"15", x"62", x"00", x"01", 
x"15", x"82", x"00", x"03", 
x"04", x"4b", x"60", x"00", 
x"08", x"63", x"ff", x"d0", 
x"04", x"42", x"18", x"00", 
x"20", x"00", x"ff", x"f7", 
x"21", x"00", x"00", x"01", 
x"10", x"40", x"10", x"00", 
x"33", x"e0", x"00", x"00", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2a", x"c5", 
x"47", x"a3", x"00", x"01", 
x"34", x"00", x"2b", x"53", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"41", x"1d", x"ff", x"ff", 
x"09", x"20", x"00", x"2e", 
x"25", x"09", x"00", x"2b", 
x"09", x"20", x"00", x"30", 
x"09", x"40", x"00", x"39", 
x"08", x"60", x"00", x"00", 
x"09", x"00", x"00", x"00", 
x"79", x"00", x"00", x"00", 
x"29", x"09", x"00", x"25", 
x"29", x"48", x"00", x"24", 
x"25", x"09", x"00", x"02", 
x"08", x"63", x"00", x"01", 
x"20", x"00", x"ff", x"fa", 
x"08", x"48", x"ff", x"d0", 
x"79", x"00", x"00", x"00", 
x"29", x"09", x"00", x"07", 
x"29", x"48", x"00", x"06", 
x"15", x"62", x"00", x"01", 
x"15", x"82", x"00", x"03", 
x"04", x"4b", x"60", x"00", 
x"09", x"08", x"ff", x"d0", 
x"04", x"42", x"40", x"00", 
x"20", x"00", x"ff", x"f7", 
x"c7", x"a2", x"ff", x"ff", 
x"47", x"a3", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"53", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"c0", x"7d", x"ff", x"ff", 
x"40", x"7d", x"ff", x"fe", 
x"09", x"00", x"00", x"04", 
x"c0", x"88", x"00", x"00", 
x"09", x"00", x"00", x"08", 
x"c0", x"a8", x"00", x"00", 
x"a8", x"44", x"00", x"02", 
x"8c", x"42", x"28", x"00", 
x"20", x"00", x"ff", x"fd", 
x"2c", x"60", x"00", x"03", 
x"08", x"63", x"ff", x"ff", 
x"8c", x"42", x"28", x"00", 
x"20", x"00", x"ff", x"fc", 
x"ac", x"03", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"33", x"e0", x"00", x"00", 
x"78", x"40", x"00", x"00", 
x"14", x"42", x"00", x"08", 
x"78", x"60", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"14", x"42", x"00", x"08", 
x"78", x"60", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"14", x"42", x"00", x"08", 
x"78", x"60", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"33", x"e0", x"00", x"00", 
x"78", x"40", x"00", x"00", 
x"14", x"42", x"00", x"08", 
x"78", x"60", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"14", x"42", x"00", x"08", 
x"78", x"60", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"14", x"42", x"00", x"08", 
x"78", x"60", x"00", x"00", 
x"04", x"42", x"18", x"00", 
x"47", x"a2", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"ff", 
x"33", x"e0", x"00", x"00", 
x"a8", x"40", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"02", 
x"09", x"00", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"09", x"20", x"00", x"0a", 
x"c0", x"69", x"00", x"00", 
x"ac", x"62", x"00", x"0a", 
x"84", x"42", x"18", x"00", 
x"c7", x"a2", x"ff", x"ff", 
x"40", x"5d", x"ff", x"ff", 
x"0d", x"40", x"4b", x"00", 
x"15", x"4a", x"00", x"10", 
x"0d", x"4a", x"00", x"00", 
x"10", x"42", x"50", x"00", 
x"21", x"00", x"00", x"01", 
x"10", x"40", x"10", x"00", 
x"33", x"e0", x"00", x"00", 
x"98", x"83", x"00", x"00", 
x"08", x"40", x"00", x"00", 
x"0d", x"60", x"00", x"80", 
x"15", x"6b", x"00", x"10", 
x"0d", x"6b", x"00", x"00", 
x"84", x"42", x"20", x"00", 
x"04", x"42", x"58", x"00", 
x"ac", x"62", x"ff", x"fd", 
x"47", x"a2", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2b", x"2e", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"40", x"7d", x"ff", x"ff", 
x"04", x"42", x"18", x"00", 
x"21", x"00", x"00", x"01", 
x"10", x"40", x"10", x"00", 
x"33", x"e0", x"00", x"00", 
x"2c", x"02", x"00", x"03", 
x"09", x"20", x"00", x"01", 
x"11", x"60", x"10", x"00", 
x"20", x"00", x"00", x"02", 
x"09", x"20", x"00", x"00", 
x"05", x"60", x"10", x"00", 
x"0d", x"00", x"00", x"80", 
x"15", x"08", x"00", x"10", 
x"0d", x"08", x"00", x"00", 
x"2d", x"0b", x"00", x"0c", 
x"0d", x"00", x"4b", x"00", 
x"15", x"08", x"00", x"10", 
x"0d", x"08", x"00", x"00", 
x"05", x"4b", x"40", x"00", 
x"47", x"aa", x"ff", x"ff", 
x"c0", x"5d", x"ff", x"ff", 
x"09", x"00", x"00", x"09", 
x"c0", x"68", x"00", x"00", 
x"84", x"42", x"18", x"00", 
x"21", x"20", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"80", x"40", x"00", x"00", 
x"09", x"00", x"00", x"0a", 
x"c0", x"68", x"00", x"00", 
x"05", x"00", x"58", x"00", 
x"05", x"20", x"00", x"00", 
x"0d", x"40", x"00", x"80", 
x"15", x"4a", x"00", x"10", 
x"0d", x"4a", x"00", x"00", 
x"11", x"60", x"50", x"00", 
x"84", x"42", x"18", x"00", 
x"05", x"08", x"58", x"00", 
x"2d", x"48", x"ff", x"fd", 
x"47", x"a2", x"ff", x"ff", 
x"c7", x"a2", x"ff", x"fe", 
x"0b", x"bd", x"ff", x"fd", 
x"47", x"bf", x"00", x"00", 
x"04", x"40", x"40", x"00", 
x"34", x"00", x"2b", x"53", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"03", 
x"c0", x"7d", x"ff", x"fe", 
x"40", x"5d", x"ff", x"ff", 
x"84", x"42", x"18", x"00", 
x"21", x"20", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"09", x"20", x"00", x"09", 
x"c0", x"a9", x"00", x"00", 
x"ac", x"45", x"00", x"13", 
x"09", x"20", x"00", x"0a", 
x"c0", x"89", x"00", x"00", 
x"ac", x"82", x"00", x"10", 
x"80", x"62", x"00", x"00", 
x"a8", x"40", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"02", 
x"09", x"00", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"84", x"42", x"20", x"00", 
x"84", x"42", x"28", x"00", 
x"21", x"00", x"00", x"01", 
x"98", x"42", x"00", x"00", 
x"09", x"20", x"00", x"06", 
x"c0", x"89", x"00", x"00", 
x"ac", x"43", x"00", x"03", 
x"84", x"a2", x"20", x"00", 
x"ac", x"65", x"00", x"01", 
x"80", x"45", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"9c", x"42", x"00", x"00", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"02", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"09", x"00", x"00", x"00", 
x"09", x"20", x"00", x"01", 
x"c0", x"69", x"00", x"00", 
x"a8", x"43", x"00", x"06", 
x"98", x"c3", x"00", x"00", 
x"84", x"42", x"30", x"00", 
x"21", x"00", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"09", x"00", x"00", x"01", 
x"09", x"20", x"00", x"02", 
x"c0", x"a9", x"00", x"00", 
x"a8", x"45", x"00", x"06", 
x"98", x"c2", x"00", x"00", 
x"84", x"43", x"30", x"00", 
x"21", x"00", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"09", x"00", x"00", x"01", 
x"09", x"20", x"00", x"03", 
x"c0", x"c9", x"00", x"00", 
x"ac", x"46", x"00", x"03", 
x"98", x"c2", x"00", x"00", 
x"84", x"45", x"30", x"00", 
x"20", x"00", x"00", x"35", 
x"8c", x"62", x"10", x"00", 
x"09", x"20", x"00", x"0d", 
x"c0", x"a9", x"00", x"00", 
x"8c", x"45", x"18", x"00", 
x"09", x"20", x"00", x"0c", 
x"c0", x"a9", x"00", x"00", 
x"84", x"42", x"28", x"00", 
x"8c", x"42", x"18", x"00", 
x"09", x"20", x"00", x"0b", 
x"c0", x"a9", x"00", x"00", 
x"84", x"42", x"28", x"00", 
x"8c", x"42", x"18", x"00", 
x"09", x"20", x"00", x"04", 
x"c0", x"a9", x"00", x"00", 
x"84", x"42", x"28", x"00", 
x"21", x"00", x"00", x"03", 
x"9c", x"42", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"9c", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"a8", x"40", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"02", 
x"09", x"00", x"00", x"01", 
x"9c", x"42", x"00", x"00", 
x"47", x"a8", x"ff", x"ff", 
x"0b", x"bd", x"ff", x"fe", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"02", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"02", 
x"41", x"1d", x"ff", x"ff", 
x"09", x"20", x"00", x"01", 
x"c0", x"69", x"00", x"00", 
x"a8", x"43", x"00", x"06", 
x"98", x"c3", x"00", x"00", 
x"84", x"42", x"30", x"00", 
x"21", x"00", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"01", 
x"09", x"00", x"00", x"01", 
x"09", x"20", x"00", x"02", 
x"c0", x"a9", x"00", x"00", 
x"a8", x"45", x"00", x"02", 
x"98", x"c2", x"00", x"00", 
x"84", x"43", x"30", x"00", 
x"09", x"20", x"00", x"03", 
x"c0", x"c9", x"00", x"00", 
x"ac", x"46", x"00", x"03", 
x"98", x"c2", x"00", x"00", 
x"84", x"45", x"30", x"00", 
x"20", x"00", x"ff", x"cb", 
x"8c", x"82", x"10", x"00", 
x"09", x"20", x"00", x"10", 
x"c0", x"a9", x"00", x"00", 
x"8c", x"65", x"20", x"00", 
x"09", x"20", x"00", x"0f", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"09", x"20", x"00", x"0e", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"8c", x"63", x"10", x"00", 
x"84", x"43", x"10", x"00", 
x"21", x"00", x"00", x"03", 
x"9c", x"42", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"9c", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"09", x"20", x"00", x"00", 
x"c0", x"69", x"00", x"00", 
x"80", x"a3", x"00", x"00", 
x"09", x"20", x"00", x"07", 
x"c0", x"89", x"00", x"00", 
x"09", x"20", x"00", x"05", 
x"c0", x"c9", x"00", x"00", 
x"a8", x"45", x"00", x"02", 
x"8c", x"a5", x"30", x"00", 
x"20", x"00", x"ff", x"fd", 
x"a8", x"43", x"00", x"05", 
x"a8", x"45", x"00", x"02", 
x"98", x"c5", x"00", x"00", 
x"84", x"42", x"30", x"00", 
x"8c", x"a5", x"20", x"00", 
x"20", x"00", x"ff", x"fa", 
x"33", x"e0", x"00", x"00", 
x"a8", x"40", x"00", x"02", 
x"09", x"00", x"00", x"00", 
x"20", x"00", x"00", x"02", 
x"09", x"00", x"00", x"01", 
x"9c", x"42", x"00", x"00", 
x"09", x"20", x"00", x"11", 
x"c0", x"c9", x"00", x"00", 
x"ac", x"c2", x"00", x"0b", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"4a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"21", x"00", x"00", x"03", 
x"9c", x"42", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"9c", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"09", x"20", x"00", x"12", 
x"c0", x"c9", x"00", x"00", 
x"ac", x"c2", x"00", x"13", 
x"09", x"20", x"00", x"04", 
x"c0", x"a9", x"00", x"00", 
x"84", x"c2", x"28", x"00", 
x"98", x"a5", x"00", x"00", 
x"84", x"e2", x"28", x"00", 
x"90", x"c6", x"00", x"00", 
x"8c", x"46", x"38", x"00", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"4a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"09", x"20", x"00", x"03", 
x"c0", x"a9", x"00", x"00", 
x"84", x"42", x"28", x"00", 
x"21", x"00", x"ff", x"eb", 
x"9c", x"42", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"90", x"42", x"00", x"00", 
x"0b", x"bd", x"ff", x"ff", 
x"47", x"bf", x"00", x"00", 
x"34", x"00", x"2c", x"4a", 
x"43", x"fd", x"00", x"00", 
x"0b", x"bd", x"00", x"01", 
x"98", x"c2", x"00", x"00", 
x"09", x"20", x"00", x"02", 
x"c0", x"49", x"00", x"00", 
x"84", x"42", x"30", x"00", 
x"21", x"00", x"ff", x"dd", 
x"9c", x"42", x"00", x"00", 
x"98", x"42", x"00", x"00", 
x"33", x"e0", x"00", x"00", 
x"8c", x"82", x"10", x"00", 
x"09", x"20", x"00", x"18", 
x"c0", x"a9", x"00", x"00", 
x"8c", x"65", x"20", x"00", 
x"09", x"20", x"00", x"17", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"09", x"20", x"00", x"16", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"09", x"20", x"00", x"15", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"09", x"20", x"00", x"14", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"09", x"20", x"00", x"13", 
x"c0", x"a9", x"00", x"00", 
x"84", x"63", x"28", x"00", 
x"8c", x"63", x"20", x"00", 
x"8c", x"63", x"10", x"00", 
x"84", x"43", x"10", x"00", 
x"33", x"e0", x"00", x"00", 
x"03", x"00", x"00", x"00", 
          
x"ff"
          );
          signal din_counter : std_logic_vector (31 downto 0) := x"00000471";
          type din_list_type is array (1137 downto 0) of std_logic_vector (7 downto 0);
          signal din_list : din_list_type := (
x"2d", x"37", x"30", x"20", 
x"20", x"33", x"35", x"20", 
x"2d", x"32", x"30", x"20", 
x"20", x"20", x"20", x"20", 
x"20", x"32", x"30", x"20", 
x"33", x"30", x"0a", x"31", 
x"20", x"35", x"30", x"20", 
x"35", x"30", x"0a", x"32", 
x"35", x"35", x"0a", x"30", 
x"20", x"31", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"32", x"30", 
x"20", x"20", x"32", x"30", 
x"20", x"20", x"36", x"35", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"32", 
x"30", x"20", x"20", x"34", 
x"35", x"20", x"20", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"31", x"32", x"38", 
x"20", x"32", x"31", x"30", 
x"20", x"20", x"20", x"30", 
x"0a", x"30", x"20", x"33", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"32", x"35", x"20", x"20", 
x"34", x"30", x"20", x"20", 
x"37", x"30", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"34", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"31", 
x"32", x"38", x"20", x"32", 
x"31", x"30", x"20", x"20", 
x"20", x"30", x"0a", x"30", 
x"20", x"33", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"33", x"30", 
x"20", x"20", x"33", x"30", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"2d", 
x"35", x"20", x"20", x"20", 
x"30", x"20", x"2d", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"31", x"32", x"38", 
x"20", x"32", x"31", x"31", 
x"20", x"20", x"20", x"30", 
x"0a", x"30", x"20", x"31", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"32", x"30", x"20", x"20", 
x"31", x"30", x"20", x"20", 
x"33", x"30", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"2d", x"31", x"30", x"20", 
x"20", x"38", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"31", 
x"32", x"38", x"20", x"32", 
x"31", x"31", x"20", x"20", 
x"20", x"30", x"0a", x"30", 
x"20", x"32", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"20", x"30", 
x"20", x"2d", x"31", x"2e", 
x"35", x"20", x"2d", x"31", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"20", 
x"30", x"20", x"20", x"35", 
x"30", x"20", x"20", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"31", x"32", x"38", 
x"20", x"32", x"31", x"31", 
x"20", x"20", x"20", x"30", 
x"0a", x"30", x"20", x"31", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"32", x"32", x"20", x"20", 
x"32", x"38", x"20", x"20", 
x"32", x"38", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"2d", x"35", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"20", 
x"20", x"30", x"20", x"32", 
x"31", x"31", x"20", x"32", 
x"31", x"31", x"0a", x"30", 
x"20", x"33", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"34", x"30", 
x"20", x"20", x"32", x"38", 
x"20", x"20", x"32", x"38", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"2d", 
x"35", x"20", x"20", x"20", 
x"30", x"20", x"20", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"20", x"20", x"30", 
x"20", x"32", x"31", x"31", 
x"20", x"32", x"31", x"31", 
x"0a", x"30", x"20", x"33", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"20", x"30", x"20", x"20", 
x"31", x"35", x"20", x"20", 
x"31", x"35", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"2d", x"35", x"20", 
x"20", x"20", x"30", x"20", 
x"2d", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"20", 
x"20", x"30", x"20", x"32", 
x"31", x"31", x"20", x"32", 
x"31", x"31", x"0a", x"30", 
x"20", x"33", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"31", x"35", 
x"20", x"20", x"32", x"35", 
x"20", x"20", x"32", x"35", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"2d", 
x"35", x"20", x"20", x"37", 
x"30", x"20", x"20", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"32", x"31", x"31", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"20", x"30", 
x"0a", x"30", x"20", x"31", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"20", x"35", x"20", x"20", 
x"31", x"31", x"20", x"20", 
x"34", x"35", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"33", x"35", x"20", 
x"20", x"34", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"32", 
x"31", x"31", x"20", x"31", 
x"32", x"38", x"20", x"20", 
x"20", x"30", x"0a", x"30", 
x"20", x"33", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"33", x"30", 
x"20", x"20", x"34", x"35", 
x"20", x"20", x"37", x"35", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"20", 
x"30", x"20", x"20", x"34", 
x"30", x"20", x"20", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"32", x"31", x"31", 
x"20", x"31", x"32", x"38", 
x"20", x"20", x"20", x"30", 
x"0a", x"30", x"20", x"31", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"32", x"35", x"20", x"20", 
x"34", x"31", x"20", x"20", 
x"37", x"30", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"20", x"35", x"20", 
x"20", x"34", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"20", 
x"20", x"30", x"20", x"20", 
x"20", x"30", x"20", x"20", 
x"20", x"30", x"0a", x"31", 
x"20", x"31", x"20", x"31", 
x"20", x"30", x"20", x"20", 
x"20", x"31", x"30", x"30", 
x"20", x"20", x"20", x"35", 
x"20", x"32", x"30", x"30", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"2d", x"33", 
x"35", x"20", x"31", x"35", 
x"30", x"20", x"20", x"31", 
x"20", x"31", x"2e", x"30", 
x"20", x"32", x"35", x"30", 
x"20", x"32", x"30", x"30", 
x"20", x"32", x"30", x"30", 
x"20", x"32", x"30", x"30", 
x"0a", x"30", x"20", x"33", 
x"20", x"31", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"32", x"35", x"20", x"20", 
x"31", x"30", x"20", x"20", 
x"31", x"30", x"20", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"2d", x"35", x"20", 
x"20", x"20", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"32", 
x"35", x"30", x"20", x"32", 
x"31", x"31", x"20", x"31", 
x"32", x"38", x"20", x"31", 
x"32", x"38", x"0a", x"30", 
x"20", x"33", x"20", x"32", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"32", x"35", 
x"20", x"20", x"32", x"30", 
x"20", x"20", x"32", x"30", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"20", 
x"30", x"20", x"20", x"37", 
x"30", x"20", x"20", x"31", 
x"20", x"30", x"2e", x"33", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"20", x"30", 
x"20", x"32", x"35", x"35", 
x"0a", x"32", x"20", x"33", 
x"20", x"31", x"20", x"30", 
x"09", x"20", x"20", x"20", 
x"32", x"30", x"20", x"20", 
x"32", x"30", x"20", x"20", 
x"32", x"30", x"20", x"20", 
x"31", x"30", x"30", x"20", 
x"20", x"34", x"30", x"20", 
x"31", x"32", x"30", x"20", 
x"20", x"31", x"20", x"31", 
x"2e", x"30", x"20", x"31", 
x"35", x"30", x"20", x"32", 
x"35", x"35", x"20", x"32", 
x"35", x"35", x"20", x"32", 
x"35", x"35", x"0a", x"30", 
x"20", x"32", x"20", x"32", 
x"20", x"30", x"20", x"20", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"2d", x"31", 
x"20", x"20", x"20", x"20", 
x"30", x"20", x"20", x"20", 
x"30", x"20", x"32", x"30", 
x"30", x"20", x"20", x"31", 
x"20", x"30", x"2e", x"32", 
x"20", x"20", x"20", x"30", 
x"20", x"32", x"35", x"35", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"20", x"30", 
x"20", x"20", x"20", x"20", 
x"20", x"0a", x"2d", x"31", 
x"0a", x"30", x"20", x"31", 
x"20", x"32", x"20", x"2d", 
x"31", x"0a", x"33", x"20", 
x"31", x"20", x"34", x"20", 
x"2d", x"31", x"0a", x"35", 
x"20", x"36", x"20", x"37", 
x"20", x"2d", x"31", x"0a", 
x"38", x"20", x"2d", x"31", 
x"0a", x"39", x"20", x"31", 
x"30", x"20", x"2d", x"31", 
x"0a", x"31", x"32", x"20", 
x"2d", x"31", x"0a", x"31", 
x"33", x"20", x"2d", x"31", 
x"0a", x"31", x"34", x"20", 
x"2d", x"31", x"0a", x"31", 
x"35", x"20", x"2d", x"31", 
x"0a", x"31", x"36", x"20", 
x"2d", x"31", x"0a", x"2d", 
x"31", x"0a", x"31", x"31", 
x"20", x"30", x"20", x"31", 
x"20", x"32", x"20", x"33", 
x"20", x"34", x"20", x"36", 
x"20", x"2d", x"31", x"0a", 
x"39", x"39", x"20", x"39", 
x"20", x"38", x"20", x"37", 
x"20", x"35", x"20", x"2d", 
x"31", x"0a", x"2d", x"31", 
x"0a", 
          
x"00"
          );

  BEGIN

  -- Component Instantiation
--          uut: TOP generic map (x"01ab") PORT MAP(
          uut: TOP generic map (wtime) PORT MAP(
            MCLK1 => clk,
            RS_RX => rs_rx,
            RS_TX => rs_tx,
            ZD => zd,
            ZA => za,
            XWA => xwa,
            XE1 => xe1,
            E2A => e2a,
            XE3 => xe3,
            XGA => xga,
            XZCKE => xzcke,
            ADVA => adva,
            XLBO => xlbo,
            ZZA => zza,
            XFT => xft,
            XZBE => xzbe,
            ZCLKMA => zclkma
            );

          sram : sram_sim port map (
            ZD => zd,
            ZA => za,
            XWA => xwa,
            XE1 => xe1,
            E2A => e2a,
            XE3 => xe3,
            XGA => xga,
            XZCKE => xzcke,
            ADVA => adva,
            XLBO => xlbo,
            ZZA => zza,
            XFT => xft,
            XZBE => xzbe,
            ZCLKMA => zclkma
        );


          recv: receiver generic map (wtime) port map (
            clk,
            receiver_in,
            receiver_out);
          send: sender generic map (wtime) port map (
            clk,
            sender_in,
            sender_out);

          receiver_in.rs_rx <= rs_tx;
          rs_rx <= sender_out.rs_tx;


  --  Test Bench Statements
     tb : PROCESS
     BEGIN
        clk <= '0';
        wait for 7.26 ns;
        clk <= '1';
        wait for 7.26 ns;
     END PROCESS tb;

     process (clk)
         variable sending : std_logic := '0';
     begin
         if rising_edge(clk) then
             if not sender_out.busy and sending = '0' then
                 if unsigned(counter) /= 0 then
                     counter <= std_logic_vector (unsigned(counter) - 1);
                     sender_in.data <= inst_list (to_integer(unsigned(counter)));
                     sender_in.go <= true;
                     sending := '1';
                 elsif unsigned(din_counter) /= 0 then
                     din_counter <= std_logic_vector (unsigned(din_counter) - 1);
                     sender_in.data <= din_list (to_integer(unsigned(din_counter)));
                     sender_in.go  <= true;
                     sending := '1';
                 else
                     sender_in.go <= false;
                     sending := '0';
                 end if;
             else
                 sender_in.go <= false;
                 sending := '0';
             end if;
         end if;
     end process;
  --  End Test Bench

  END;
